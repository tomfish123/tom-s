//////////////////////////////////////////////////////////////////////////////////
// Description:
//////////////////////////////////////////////////////////////////////////////////

module pdec_rom_depth
#(parameter D=16384,
  parameter W=32,
  parameter RD_TYPE=0) //0=delay address by 1T;1=delay rdata
(
  input                 clk,
  input                 ce,   //high active
  input                 we,   //high active
  input  [$clog2(D)-1:0]addr,
  input  [W-1:0]        wdata,
  output [W-1:0]        rdata
);

  wire [W-1:0] mem[0:D-1];
  //----initial
  assign mem[0   ] = 4'h0; 
  assign mem[1   ] = 4'h1;
  assign mem[2   ] = 4'h0;
  assign mem[3   ] = 4'h2;
  assign mem[4   ] = 4'h0;
  assign mem[5   ] = 4'h1;
  assign mem[6   ] = 4'h0;
  assign mem[7   ] = 4'h3;
  assign mem[8   ] = 4'h0;
  assign mem[9   ] = 4'h1;
  assign mem[10  ] = 4'h0;
  assign mem[11  ] = 4'h2;
  assign mem[12  ] = 4'h0;
  assign mem[13  ] = 4'h1;
  assign mem[14  ] = 4'h0;
  assign mem[15  ] = 4'h4;
  assign mem[16  ] = 4'h0;
  assign mem[17  ] = 4'h1;
  assign mem[18  ] = 4'h0;
  assign mem[19  ] = 4'h2;
  assign mem[20  ] = 4'h0;
  assign mem[21  ] = 4'h1;
  assign mem[22  ] = 4'h0;
  assign mem[23  ] = 4'h3;
  assign mem[24  ] = 4'h0;
  assign mem[25  ] = 4'h1;
  assign mem[26  ] = 4'h0;
  assign mem[27  ] = 4'h2;
  assign mem[28  ] = 4'h0;
  assign mem[29  ] = 4'h1;
  assign mem[30  ] = 4'h0;
  assign mem[31  ] = 4'h5;
  assign mem[32  ] = 4'h0;
  assign mem[33  ] = 4'h1;
  assign mem[34  ] = 4'h0;
  assign mem[35  ] = 4'h2;
  assign mem[36  ] = 4'h0;
  assign mem[37  ] = 4'h1;
  assign mem[38  ] = 4'h0;
  assign mem[39  ] = 4'h3;
  assign mem[40  ] = 4'h0;
  assign mem[41  ] = 4'h1;
  assign mem[42  ] = 4'h0;
  assign mem[43  ] = 4'h2;
  assign mem[44  ] = 4'h0;
  assign mem[45  ] = 4'h1;
  assign mem[46  ] = 4'h0;
  assign mem[47  ] = 4'h4;
  assign mem[48  ] = 4'h0;
  assign mem[49  ] = 4'h1;
  assign mem[50  ] = 4'h0;
  assign mem[51  ] = 4'h2;
  assign mem[52  ] = 4'h0;
  assign mem[53  ] = 4'h1;
  assign mem[54  ] = 4'h0;
  assign mem[55  ] = 4'h3;
  assign mem[56  ] = 4'h0;
  assign mem[57  ] = 4'h1;
  assign mem[58  ] = 4'h0;
  assign mem[59  ] = 4'h2;
  assign mem[60  ] = 4'h0;
  assign mem[61  ] = 4'h1;
  assign mem[62  ] = 4'h0;
  assign mem[63  ] = 4'h6;
  assign mem[64  ] = 4'h0;
  assign mem[65  ] = 4'h1;
  assign mem[66  ] = 4'h0;
  assign mem[67  ] = 4'h2;
  assign mem[68  ] = 4'h0;
  assign mem[69  ] = 4'h1;
  assign mem[70  ] = 4'h0;
  assign mem[71  ] = 4'h3;
  assign mem[72  ] = 4'h0;
  assign mem[73  ] = 4'h1;
  assign mem[74  ] = 4'h0;
  assign mem[75  ] = 4'h2;
  assign mem[76  ] = 4'h0;
  assign mem[77  ] = 4'h1;
  assign mem[78  ] = 4'h0;
  assign mem[79  ] = 4'h4;
  assign mem[80  ] = 4'h0;
  assign mem[81  ] = 4'h1;
  assign mem[82  ] = 4'h0;
  assign mem[83  ] = 4'h2;
  assign mem[84  ] = 4'h0;
  assign mem[85  ] = 4'h1;
  assign mem[86  ] = 4'h0;
  assign mem[87  ] = 4'h3;
  assign mem[88  ] = 4'h0;
  assign mem[89  ] = 4'h1;
  assign mem[90  ] = 4'h0;
  assign mem[91  ] = 4'h2;
  assign mem[92  ] = 4'h0;
  assign mem[93  ] = 4'h1;
  assign mem[94  ] = 4'h0;
  assign mem[95  ] = 4'h5;
  assign mem[96  ] = 4'h0;
  assign mem[97  ] = 4'h1;
  assign mem[98  ] = 4'h0;
  assign mem[99  ] = 4'h2;
  assign mem[100 ] = 4'h0;
  assign mem[101 ] = 4'h1;
  assign mem[102 ] = 4'h0;
  assign mem[103 ] = 4'h3;
  assign mem[104 ] = 4'h0;
  assign mem[105 ] = 4'h1;
  assign mem[106 ] = 4'h0;
  assign mem[107 ] = 4'h2;
  assign mem[108 ] = 4'h0;
  assign mem[109 ] = 4'h1;
  assign mem[110 ] = 4'h0;
  assign mem[111 ] = 4'h4;
  assign mem[112 ] = 4'h0;
  assign mem[113 ] = 4'h1;
  assign mem[114 ] = 4'h0;
  assign mem[115 ] = 4'h2;
  assign mem[116 ] = 4'h0;
  assign mem[117 ] = 4'h1;
  assign mem[118 ] = 4'h0;
  assign mem[119 ] = 4'h3;
  assign mem[120 ] = 4'h0;
  assign mem[121 ] = 4'h1;
  assign mem[122 ] = 4'h0;
  assign mem[123 ] = 4'h2;
  assign mem[124 ] = 4'h0;
  assign mem[125 ] = 4'h1;
  assign mem[126 ] = 4'h0;
  assign mem[127 ] = 4'h7;
  assign mem[128 ] = 4'h0;
  assign mem[129 ] = 4'h1;
  assign mem[130 ] = 4'h0;
  assign mem[131 ] = 4'h2;
  assign mem[132 ] = 4'h0;
  assign mem[133 ] = 4'h1;
  assign mem[134 ] = 4'h0;
  assign mem[135 ] = 4'h3;
  assign mem[136 ] = 4'h0;
  assign mem[137 ] = 4'h1;
  assign mem[138 ] = 4'h0;
  assign mem[139 ] = 4'h2;
  assign mem[140 ] = 4'h0;
  assign mem[141 ] = 4'h1;
  assign mem[142 ] = 4'h0;
  assign mem[143 ] = 4'h4;
  assign mem[144 ] = 4'h0;
  assign mem[145 ] = 4'h1;
  assign mem[146 ] = 4'h0;
  assign mem[147 ] = 4'h2;
  assign mem[148 ] = 4'h0;
  assign mem[149 ] = 4'h1;
  assign mem[150 ] = 4'h0;
  assign mem[151 ] = 4'h3;
  assign mem[152 ] = 4'h0;
  assign mem[153 ] = 4'h1;
  assign mem[154 ] = 4'h0;
  assign mem[155 ] = 4'h2;
  assign mem[156 ] = 4'h0;
  assign mem[157 ] = 4'h1;
  assign mem[158 ] = 4'h0;
  assign mem[159 ] = 4'h5;
  assign mem[160 ] = 4'h0;
  assign mem[161 ] = 4'h1;
  assign mem[162 ] = 4'h0;
  assign mem[163 ] = 4'h2;
  assign mem[164 ] = 4'h0;
  assign mem[165 ] = 4'h1;
  assign mem[166 ] = 4'h0;
  assign mem[167 ] = 4'h3;
  assign mem[168 ] = 4'h0;
  assign mem[169 ] = 4'h1;
  assign mem[170 ] = 4'h0;
  assign mem[171 ] = 4'h2;
  assign mem[172 ] = 4'h0;
  assign mem[173 ] = 4'h1;
  assign mem[174 ] = 4'h0;
  assign mem[175 ] = 4'h4;
  assign mem[176 ] = 4'h0;
  assign mem[177 ] = 4'h1;
  assign mem[178 ] = 4'h0;
  assign mem[179 ] = 4'h2;
  assign mem[180 ] = 4'h0;
  assign mem[181 ] = 4'h1;
  assign mem[182 ] = 4'h0;
  assign mem[183 ] = 4'h3;
  assign mem[184 ] = 4'h0;
  assign mem[185 ] = 4'h1;
  assign mem[186 ] = 4'h0;
  assign mem[187 ] = 4'h2;
  assign mem[188 ] = 4'h0;
  assign mem[189 ] = 4'h1;
  assign mem[190 ] = 4'h0;
  assign mem[191 ] = 4'h6;
  assign mem[192 ] = 4'h0;
  assign mem[193 ] = 4'h1;
  assign mem[194 ] = 4'h0;
  assign mem[195 ] = 4'h2;
  assign mem[196 ] = 4'h0;
  assign mem[197 ] = 4'h1;
  assign mem[198 ] = 4'h0;
  assign mem[199 ] = 4'h3;
  assign mem[200 ] = 4'h0;
  assign mem[201 ] = 4'h1;
  assign mem[202 ] = 4'h0;
  assign mem[203 ] = 4'h2;
  assign mem[204 ] = 4'h0;
  assign mem[205 ] = 4'h1;
  assign mem[206 ] = 4'h0;
  assign mem[207 ] = 4'h4;
  assign mem[208 ] = 4'h0;
  assign mem[209 ] = 4'h1;
  assign mem[210 ] = 4'h0;
  assign mem[211 ] = 4'h2;
  assign mem[212 ] = 4'h0;
  assign mem[213 ] = 4'h1;
  assign mem[214 ] = 4'h0;
  assign mem[215 ] = 4'h3;
  assign mem[216 ] = 4'h0;
  assign mem[217 ] = 4'h1;
  assign mem[218 ] = 4'h0;
  assign mem[219 ] = 4'h2;
  assign mem[220 ] = 4'h0;
  assign mem[221 ] = 4'h1;
  assign mem[222 ] = 4'h0;
  assign mem[223 ] = 4'h5;
  assign mem[224 ] = 4'h0;
  assign mem[225 ] = 4'h1;
  assign mem[226 ] = 4'h0;
  assign mem[227 ] = 4'h2;
  assign mem[228 ] = 4'h0;
  assign mem[229 ] = 4'h1;
  assign mem[230 ] = 4'h0;
  assign mem[231 ] = 4'h3;
  assign mem[232 ] = 4'h0;
  assign mem[233 ] = 4'h1;
  assign mem[234 ] = 4'h0;
  assign mem[235 ] = 4'h2;
  assign mem[236 ] = 4'h0;
  assign mem[237 ] = 4'h1;
  assign mem[238 ] = 4'h0;
  assign mem[239 ] = 4'h4;
  assign mem[240 ] = 4'h0;
  assign mem[241 ] = 4'h1;
  assign mem[242 ] = 4'h0;
  assign mem[243 ] = 4'h2;
  assign mem[244 ] = 4'h0;
  assign mem[245 ] = 4'h1;
  assign mem[246 ] = 4'h0;
  assign mem[247 ] = 4'h3;
  assign mem[248 ] = 4'h0;
  assign mem[249 ] = 4'h1;
  assign mem[250 ] = 4'h0;
  assign mem[251 ] = 4'h2;
  assign mem[252 ] = 4'h0;
  assign mem[253 ] = 4'h1;
  assign mem[254 ] = 4'h0;
  assign mem[255 ] = 4'h8;
  assign mem[256 ] = 4'h0;
  assign mem[257 ] = 4'h1;
  assign mem[258 ] = 4'h0;
  assign mem[259 ] = 4'h2;
  assign mem[260 ] = 4'h0;
  assign mem[261 ] = 4'h1;
  assign mem[262 ] = 4'h0;
  assign mem[263 ] = 4'h3;
  assign mem[264 ] = 4'h0;
  assign mem[265 ] = 4'h1;
  assign mem[266 ] = 4'h0;
  assign mem[267 ] = 4'h2;
  assign mem[268 ] = 4'h0;
  assign mem[269 ] = 4'h1;
  assign mem[270 ] = 4'h0;
  assign mem[271 ] = 4'h4;
  assign mem[272 ] = 4'h0;
  assign mem[273 ] = 4'h1;
  assign mem[274 ] = 4'h0;
  assign mem[275 ] = 4'h2;
  assign mem[276 ] = 4'h0;
  assign mem[277 ] = 4'h1;
  assign mem[278 ] = 4'h0;
  assign mem[279 ] = 4'h3;
  assign mem[280 ] = 4'h0;
  assign mem[281 ] = 4'h1;
  assign mem[282 ] = 4'h0;
  assign mem[283 ] = 4'h2;
  assign mem[284 ] = 4'h0;
  assign mem[285 ] = 4'h1;
  assign mem[286 ] = 4'h0;
  assign mem[287 ] = 4'h5;
  assign mem[288 ] = 4'h0;
  assign mem[289 ] = 4'h1;
  assign mem[290 ] = 4'h0;
  assign mem[291 ] = 4'h2;
  assign mem[292 ] = 4'h0;
  assign mem[293 ] = 4'h1;
  assign mem[294 ] = 4'h0;
  assign mem[295 ] = 4'h3;
  assign mem[296 ] = 4'h0;
  assign mem[297 ] = 4'h1;
  assign mem[298 ] = 4'h0;
  assign mem[299 ] = 4'h2;
  assign mem[300 ] = 4'h0;
  assign mem[301 ] = 4'h1;
  assign mem[302 ] = 4'h0;
  assign mem[303 ] = 4'h4;
  assign mem[304 ] = 4'h0;
  assign mem[305 ] = 4'h1;
  assign mem[306 ] = 4'h0;
  assign mem[307 ] = 4'h2;
  assign mem[308 ] = 4'h0;
  assign mem[309 ] = 4'h1;
  assign mem[310 ] = 4'h0;
  assign mem[311 ] = 4'h3;
  assign mem[312 ] = 4'h0;
  assign mem[313 ] = 4'h1;
  assign mem[314 ] = 4'h0;
  assign mem[315 ] = 4'h2;
  assign mem[316 ] = 4'h0;
  assign mem[317 ] = 4'h1;
  assign mem[318 ] = 4'h0;
  assign mem[319 ] = 4'h6;
  assign mem[320 ] = 4'h0;
  assign mem[321 ] = 4'h1;
  assign mem[322 ] = 4'h0;
  assign mem[323 ] = 4'h2;
  assign mem[324 ] = 4'h0;
  assign mem[325 ] = 4'h1;
  assign mem[326 ] = 4'h0;
  assign mem[327 ] = 4'h3;
  assign mem[328 ] = 4'h0;
  assign mem[329 ] = 4'h1;
  assign mem[330 ] = 4'h0;
  assign mem[331 ] = 4'h2;
  assign mem[332 ] = 4'h0;
  assign mem[333 ] = 4'h1;
  assign mem[334 ] = 4'h0;
  assign mem[335 ] = 4'h4;
  assign mem[336 ] = 4'h0;
  assign mem[337 ] = 4'h1;
  assign mem[338 ] = 4'h0;
  assign mem[339 ] = 4'h2;
  assign mem[340 ] = 4'h0;
  assign mem[341 ] = 4'h1;
  assign mem[342 ] = 4'h0;
  assign mem[343 ] = 4'h3;
  assign mem[344 ] = 4'h0;
  assign mem[345 ] = 4'h1;
  assign mem[346 ] = 4'h0;
  assign mem[347 ] = 4'h2;
  assign mem[348 ] = 4'h0;
  assign mem[349 ] = 4'h1;
  assign mem[350 ] = 4'h0;
  assign mem[351 ] = 4'h5;
  assign mem[352 ] = 4'h0;
  assign mem[353 ] = 4'h1;
  assign mem[354 ] = 4'h0;
  assign mem[355 ] = 4'h2;
  assign mem[356 ] = 4'h0;
  assign mem[357 ] = 4'h1;
  assign mem[358 ] = 4'h0;
  assign mem[359 ] = 4'h3;
  assign mem[360 ] = 4'h0;
  assign mem[361 ] = 4'h1;
  assign mem[362 ] = 4'h0;
  assign mem[363 ] = 4'h2;
  assign mem[364 ] = 4'h0;
  assign mem[365 ] = 4'h1;
  assign mem[366 ] = 4'h0;
  assign mem[367 ] = 4'h4;
  assign mem[368 ] = 4'h0;
  assign mem[369 ] = 4'h1;
  assign mem[370 ] = 4'h0;
  assign mem[371 ] = 4'h2;
  assign mem[372 ] = 4'h0;
  assign mem[373 ] = 4'h1;
  assign mem[374 ] = 4'h0;
  assign mem[375 ] = 4'h3;
  assign mem[376 ] = 4'h0;
  assign mem[377 ] = 4'h1;
  assign mem[378 ] = 4'h0;
  assign mem[379 ] = 4'h2;
  assign mem[380 ] = 4'h0;
  assign mem[381 ] = 4'h1;
  assign mem[382 ] = 4'h0;
  assign mem[383 ] = 4'h7;
  assign mem[384 ] = 4'h0;
  assign mem[385 ] = 4'h1;
  assign mem[386 ] = 4'h0;
  assign mem[387 ] = 4'h2;
  assign mem[388 ] = 4'h0;
  assign mem[389 ] = 4'h1;
  assign mem[390 ] = 4'h0;
  assign mem[391 ] = 4'h3;
  assign mem[392 ] = 4'h0;
  assign mem[393 ] = 4'h1;
  assign mem[394 ] = 4'h0;
  assign mem[395 ] = 4'h2;
  assign mem[396 ] = 4'h0;
  assign mem[397 ] = 4'h1;
  assign mem[398 ] = 4'h0;
  assign mem[399 ] = 4'h4;
  assign mem[400 ] = 4'h0;
  assign mem[401 ] = 4'h1;
  assign mem[402 ] = 4'h0;
  assign mem[403 ] = 4'h2;
  assign mem[404 ] = 4'h0;
  assign mem[405 ] = 4'h1;
  assign mem[406 ] = 4'h0;
  assign mem[407 ] = 4'h3;
  assign mem[408 ] = 4'h0;
  assign mem[409 ] = 4'h1;
  assign mem[410 ] = 4'h0;
  assign mem[411 ] = 4'h2;
  assign mem[412 ] = 4'h0;
  assign mem[413 ] = 4'h1;
  assign mem[414 ] = 4'h0;
  assign mem[415 ] = 4'h5;
  assign mem[416 ] = 4'h0;
  assign mem[417 ] = 4'h1;
  assign mem[418 ] = 4'h0;
  assign mem[419 ] = 4'h2;
  assign mem[420 ] = 4'h0;
  assign mem[421 ] = 4'h1;
  assign mem[422 ] = 4'h0;
  assign mem[423 ] = 4'h3;
  assign mem[424 ] = 4'h0;
  assign mem[425 ] = 4'h1;
  assign mem[426 ] = 4'h0;
  assign mem[427 ] = 4'h2;
  assign mem[428 ] = 4'h0;
  assign mem[429 ] = 4'h1;
  assign mem[430 ] = 4'h0;
  assign mem[431 ] = 4'h4;
  assign mem[432 ] = 4'h0;
  assign mem[433 ] = 4'h1;
  assign mem[434 ] = 4'h0;
  assign mem[435 ] = 4'h2;
  assign mem[436 ] = 4'h0;
  assign mem[437 ] = 4'h1;
  assign mem[438 ] = 4'h0;
  assign mem[439 ] = 4'h3;
  assign mem[440 ] = 4'h0;
  assign mem[441 ] = 4'h1;
  assign mem[442 ] = 4'h0;
  assign mem[443 ] = 4'h2;
  assign mem[444 ] = 4'h0;
  assign mem[445 ] = 4'h1;
  assign mem[446 ] = 4'h0;
  assign mem[447 ] = 4'h6;
  assign mem[448 ] = 4'h0;
  assign mem[449 ] = 4'h1;
  assign mem[450 ] = 4'h0;
  assign mem[451 ] = 4'h2;
  assign mem[452 ] = 4'h0;
  assign mem[453 ] = 4'h1;
  assign mem[454 ] = 4'h0;
  assign mem[455 ] = 4'h3;
  assign mem[456 ] = 4'h0;
  assign mem[457 ] = 4'h1;
  assign mem[458 ] = 4'h0;
  assign mem[459 ] = 4'h2;
  assign mem[460 ] = 4'h0;
  assign mem[461 ] = 4'h1;
  assign mem[462 ] = 4'h0;
  assign mem[463 ] = 4'h4;
  assign mem[464 ] = 4'h0;
  assign mem[465 ] = 4'h1;
  assign mem[466 ] = 4'h0;
  assign mem[467 ] = 4'h2;
  assign mem[468 ] = 4'h0;
  assign mem[469 ] = 4'h1;
  assign mem[470 ] = 4'h0;
  assign mem[471 ] = 4'h3;
  assign mem[472 ] = 4'h0;
  assign mem[473 ] = 4'h1;
  assign mem[474 ] = 4'h0;
  assign mem[475 ] = 4'h2;
  assign mem[476 ] = 4'h0;
  assign mem[477 ] = 4'h1;
  assign mem[478 ] = 4'h0;
  assign mem[479 ] = 4'h5;
  assign mem[480 ] = 4'h0;
  assign mem[481 ] = 4'h1;
  assign mem[482 ] = 4'h0;
  assign mem[483 ] = 4'h2;
  assign mem[484 ] = 4'h0;
  assign mem[485 ] = 4'h1;
  assign mem[486 ] = 4'h0;
  assign mem[487 ] = 4'h3;
  assign mem[488 ] = 4'h0;
  assign mem[489 ] = 4'h1;
  assign mem[490 ] = 4'h0;
  assign mem[491 ] = 4'h2;
  assign mem[492 ] = 4'h0;
  assign mem[493 ] = 4'h1;
  assign mem[494 ] = 4'h0;
  assign mem[495 ] = 4'h4;
  assign mem[496 ] = 4'h0;
  assign mem[497 ] = 4'h1;
  assign mem[498 ] = 4'h0;
  assign mem[499 ] = 4'h2;
  assign mem[500 ] = 4'h0;
  assign mem[501 ] = 4'h1;
  assign mem[502 ] = 4'h0;
  assign mem[503 ] = 4'h3;
  assign mem[504 ] = 4'h0;
  assign mem[505 ] = 4'h1;
  assign mem[506 ] = 4'h0;
  assign mem[507 ] = 4'h2;
  assign mem[508 ] = 4'h0;
  assign mem[509 ] = 4'h1;
  assign mem[510 ] = 4'h0;
  assign mem[511 ] = 4'h0;
  //----
  generate 
  if (RD_TYPE==0)
  begin:U_type0
    reg [$clog2(D)-1:0]addr_d1;

    always @(posedge clk)
    begin
      if((!we) & ce)
        addr_d1 <= addr;
    end

    assign rdata = mem[addr_d1];
  end
  else 
  begin:U_type1

    reg [W-1:0]rdata_int;
    always @(posedge clk)
    begin
      if((!we) & ce)
        rdata_int <= mem[addr];
    end

    assign rdata = rdata_int;
  end
  endgenerate
endmodule
