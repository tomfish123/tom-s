//////////////////////////////////////////////////////////////////////////////////
// Description:
//////////////////////////////////////////////////////////////////////////////////

module pdec_rom_stage_bd
#(parameter D=16384,
  parameter W=32,
  parameter RD_TYPE=0) //0=delay address by 1T;1=delay rdata
(
  input                 clk,
  input                 ce,   //high active
  input                 we,   //high active
  input  [$clog2(D)-1:0]addr,
  input  [W-1:0]        wdata,
  output [W-1:0]        rdata
);

  wire [W-1:0] mem[0:D-1]/*synthesis syn_ramstyle="block_ram" */;
  //----intial
  assign mem[0   ] = 5'h1b; 
  assign mem[1   ] = 5'h1a;
  assign mem[2   ] = 5'h19;
  assign mem[3   ] = 5'h18;
  assign mem[4   ] = 5'h17;
  assign mem[5   ] = 5'h16;
  assign mem[6   ] = 5'h15;
  assign mem[7   ] = 5'h14;
  assign mem[8   ] = 5'h13;
  assign mem[9   ] = 5'h12;
  assign mem[10  ] = 5'h11;
  assign mem[11  ] = 5'h10;
  assign mem[12  ] = 5'h00;
  assign mem[13  ] = 5'h01;
  assign mem[14  ] = 5'h10;
  assign mem[15  ] = 5'h00;
  assign mem[16  ] = 5'h02;
  assign mem[17  ] = 5'h11;
  assign mem[18  ] = 5'h10;
  assign mem[19  ] = 5'h00;
  assign mem[20  ] = 5'h01;
  assign mem[21  ] = 5'h10;
  assign mem[22  ] = 5'h00;
  assign mem[23  ] = 5'h03;
  assign mem[24  ] = 5'h12;
  assign mem[25  ] = 5'h11;
  assign mem[26  ] = 5'h10;
  assign mem[27  ] = 5'h00;
  assign mem[28  ] = 5'h01;
  assign mem[29  ] = 5'h10;
  assign mem[30  ] = 5'h00;
  assign mem[31  ] = 5'h02;
  assign mem[32  ] = 5'h11;
  assign mem[33  ] = 5'h10;
  assign mem[34  ] = 5'h00;
  assign mem[35  ] = 5'h01;
  assign mem[36  ] = 5'h10;
  assign mem[37  ] = 5'h00;
  assign mem[38  ] = 5'h04;
  assign mem[39  ] = 5'h13;
  assign mem[40  ] = 5'h12;
  assign mem[41  ] = 5'h11;
  assign mem[42  ] = 5'h10;
  assign mem[43  ] = 5'h00;
  assign mem[44  ] = 5'h01;
  assign mem[45  ] = 5'h10;
  assign mem[46  ] = 5'h00;
  assign mem[47  ] = 5'h02;
  assign mem[48  ] = 5'h11;
  assign mem[49  ] = 5'h10;
  assign mem[50  ] = 5'h00;
  assign mem[51  ] = 5'h01;
  assign mem[52  ] = 5'h10;
  assign mem[53  ] = 5'h00;
  assign mem[54  ] = 5'h03;
  assign mem[55  ] = 5'h12;
  assign mem[56  ] = 5'h11;
  assign mem[57  ] = 5'h10;
  assign mem[58  ] = 5'h00;
  assign mem[59  ] = 5'h01;
  assign mem[60  ] = 5'h10;
  assign mem[61  ] = 5'h00;
  assign mem[62  ] = 5'h02;
  assign mem[63  ] = 5'h11;
  assign mem[64  ] = 5'h10;
  assign mem[65  ] = 5'h00;
  assign mem[66  ] = 5'h01;
  assign mem[67  ] = 5'h10;
  assign mem[68  ] = 5'h00;
  assign mem[69  ] = 5'h05;
  assign mem[70  ] = 5'h14;
  assign mem[71  ] = 5'h13;
  assign mem[72  ] = 5'h12;
  assign mem[73  ] = 5'h11;
  assign mem[74  ] = 5'h10;
  assign mem[75  ] = 5'h00;
  assign mem[76  ] = 5'h01;
  assign mem[77  ] = 5'h10;
  assign mem[78  ] = 5'h00;
  assign mem[79  ] = 5'h02;
  assign mem[80  ] = 5'h11;
  assign mem[81  ] = 5'h10;
  assign mem[82  ] = 5'h00;
  assign mem[83  ] = 5'h01;
  assign mem[84  ] = 5'h10;
  assign mem[85  ] = 5'h00;
  assign mem[86  ] = 5'h03;
  assign mem[87  ] = 5'h12;
  assign mem[88  ] = 5'h11;
  assign mem[89  ] = 5'h10;
  assign mem[90  ] = 5'h00;
  assign mem[91  ] = 5'h01;
  assign mem[92  ] = 5'h10;
  assign mem[93  ] = 5'h00;
  assign mem[94  ] = 5'h02;
  assign mem[95  ] = 5'h11;
  assign mem[96  ] = 5'h10;
  assign mem[97  ] = 5'h00;
  assign mem[98  ] = 5'h01;
  assign mem[99  ] = 5'h10;
  assign mem[100 ] = 5'h00;
  assign mem[101 ] = 5'h04;
  assign mem[102 ] = 5'h13;
  assign mem[103 ] = 5'h12;
  assign mem[104 ] = 5'h11;
  assign mem[105 ] = 5'h10;
  assign mem[106 ] = 5'h00;
  assign mem[107 ] = 5'h01;
  assign mem[108 ] = 5'h10;
  assign mem[109 ] = 5'h00;
  assign mem[110 ] = 5'h02;
  assign mem[111 ] = 5'h11;
  assign mem[112 ] = 5'h10;
  assign mem[113 ] = 5'h00;
  assign mem[114 ] = 5'h01;
  assign mem[115 ] = 5'h10;
  assign mem[116 ] = 5'h00;
  assign mem[117 ] = 5'h03;
  assign mem[118 ] = 5'h12;
  assign mem[119 ] = 5'h11;
  assign mem[120 ] = 5'h10;
  assign mem[121 ] = 5'h00;
  assign mem[122 ] = 5'h01;
  assign mem[123 ] = 5'h10;
  assign mem[124 ] = 5'h00;
  assign mem[125 ] = 5'h02;
  assign mem[126 ] = 5'h11;
  assign mem[127 ] = 5'h10;
  assign mem[128 ] = 5'h00;
  assign mem[129 ] = 5'h01;
  assign mem[130 ] = 5'h10;
  assign mem[131 ] = 5'h00;
  assign mem[132 ] = 5'h06;
  assign mem[133 ] = 5'h15;
  assign mem[134 ] = 5'h14;
  assign mem[135 ] = 5'h13;
  assign mem[136 ] = 5'h12;
  assign mem[137 ] = 5'h11;
  assign mem[138 ] = 5'h10;
  assign mem[139 ] = 5'h00;
  assign mem[140 ] = 5'h01;
  assign mem[141 ] = 5'h10;
  assign mem[142 ] = 5'h00;
  assign mem[143 ] = 5'h02;
  assign mem[144 ] = 5'h11;
  assign mem[145 ] = 5'h10;
  assign mem[146 ] = 5'h00;
  assign mem[147 ] = 5'h01;
  assign mem[148 ] = 5'h10;
  assign mem[149 ] = 5'h00;
  assign mem[150 ] = 5'h03;
  assign mem[151 ] = 5'h12;
  assign mem[152 ] = 5'h11;
  assign mem[153 ] = 5'h10;
  assign mem[154 ] = 5'h00;
  assign mem[155 ] = 5'h01;
  assign mem[156 ] = 5'h10;
  assign mem[157 ] = 5'h00;
  assign mem[158 ] = 5'h02;
  assign mem[159 ] = 5'h11;
  assign mem[160 ] = 5'h10;
  assign mem[161 ] = 5'h00;
  assign mem[162 ] = 5'h01;
  assign mem[163 ] = 5'h10;
  assign mem[164 ] = 5'h00;
  assign mem[165 ] = 5'h04;
  assign mem[166 ] = 5'h13;
  assign mem[167 ] = 5'h12;
  assign mem[168 ] = 5'h11;
  assign mem[169 ] = 5'h10;
  assign mem[170 ] = 5'h00;
  assign mem[171 ] = 5'h01;
  assign mem[172 ] = 5'h10;
  assign mem[173 ] = 5'h00;
  assign mem[174 ] = 5'h02;
  assign mem[175 ] = 5'h11;
  assign mem[176 ] = 5'h10;
  assign mem[177 ] = 5'h00;
  assign mem[178 ] = 5'h01;
  assign mem[179 ] = 5'h10;
  assign mem[180 ] = 5'h00;
  assign mem[181 ] = 5'h03;
  assign mem[182 ] = 5'h12;
  assign mem[183 ] = 5'h11;
  assign mem[184 ] = 5'h10;
  assign mem[185 ] = 5'h00;
  assign mem[186 ] = 5'h01;
  assign mem[187 ] = 5'h10;
  assign mem[188 ] = 5'h00;
  assign mem[189 ] = 5'h02;
  assign mem[190 ] = 5'h11;
  assign mem[191 ] = 5'h10;
  assign mem[192 ] = 5'h00;
  assign mem[193 ] = 5'h01;
  assign mem[194 ] = 5'h10;
  assign mem[195 ] = 5'h00;
  assign mem[196 ] = 5'h05;
  assign mem[197 ] = 5'h14;
  assign mem[198 ] = 5'h13;
  assign mem[199 ] = 5'h12;
  assign mem[200 ] = 5'h11;
  assign mem[201 ] = 5'h10;
  assign mem[202 ] = 5'h00;
  assign mem[203 ] = 5'h01;
  assign mem[204 ] = 5'h10;
  assign mem[205 ] = 5'h00;
  assign mem[206 ] = 5'h02;
  assign mem[207 ] = 5'h11;
  assign mem[208 ] = 5'h10;
  assign mem[209 ] = 5'h00;
  assign mem[210 ] = 5'h01;
  assign mem[211 ] = 5'h10;
  assign mem[212 ] = 5'h00;
  assign mem[213 ] = 5'h03;
  assign mem[214 ] = 5'h12;
  assign mem[215 ] = 5'h11;
  assign mem[216 ] = 5'h10;
  assign mem[217 ] = 5'h00;
  assign mem[218 ] = 5'h01;
  assign mem[219 ] = 5'h10;
  assign mem[220 ] = 5'h00;
  assign mem[221 ] = 5'h02;
  assign mem[222 ] = 5'h11;
  assign mem[223 ] = 5'h10;
  assign mem[224 ] = 5'h00;
  assign mem[225 ] = 5'h01;
  assign mem[226 ] = 5'h10;
  assign mem[227 ] = 5'h00;
  assign mem[228 ] = 5'h04;
  assign mem[229 ] = 5'h13;
  assign mem[230 ] = 5'h12;
  assign mem[231 ] = 5'h11;
  assign mem[232 ] = 5'h10;
  assign mem[233 ] = 5'h00;
  assign mem[234 ] = 5'h01;
  assign mem[235 ] = 5'h10;
  assign mem[236 ] = 5'h00;
  assign mem[237 ] = 5'h02;
  assign mem[238 ] = 5'h11;
  assign mem[239 ] = 5'h10;
  assign mem[240 ] = 5'h00;
  assign mem[241 ] = 5'h01;
  assign mem[242 ] = 5'h10;
  assign mem[243 ] = 5'h00;
  assign mem[244 ] = 5'h03;
  assign mem[245 ] = 5'h12;
  assign mem[246 ] = 5'h11;
  assign mem[247 ] = 5'h10;
  assign mem[248 ] = 5'h00;
  assign mem[249 ] = 5'h01;
  assign mem[250 ] = 5'h10;
  assign mem[251 ] = 5'h00;
  assign mem[252 ] = 5'h02;
  assign mem[253 ] = 5'h11;
  assign mem[254 ] = 5'h10;
  assign mem[255 ] = 5'h00;
  assign mem[256 ] = 5'h01;
  assign mem[257 ] = 5'h10;
  assign mem[258 ] = 5'h00;
  assign mem[259 ] = 5'h07;
  assign mem[260 ] = 5'h16;
  assign mem[261 ] = 5'h15;
  assign mem[262 ] = 5'h14;
  assign mem[263 ] = 5'h13;
  assign mem[264 ] = 5'h12;
  assign mem[265 ] = 5'h11;
  assign mem[266 ] = 5'h10;
  assign mem[267 ] = 5'h00;
  assign mem[268 ] = 5'h01;
  assign mem[269 ] = 5'h10;
  assign mem[270 ] = 5'h00;
  assign mem[271 ] = 5'h02;
  assign mem[272 ] = 5'h11;
  assign mem[273 ] = 5'h10;
  assign mem[274 ] = 5'h00;
  assign mem[275 ] = 5'h01;
  assign mem[276 ] = 5'h10;
  assign mem[277 ] = 5'h00;
  assign mem[278 ] = 5'h03;
  assign mem[279 ] = 5'h12;
  assign mem[280 ] = 5'h11;
  assign mem[281 ] = 5'h10;
  assign mem[282 ] = 5'h00;
  assign mem[283 ] = 5'h01;
  assign mem[284 ] = 5'h10;
  assign mem[285 ] = 5'h00;
  assign mem[286 ] = 5'h02;
  assign mem[287 ] = 5'h11;
  assign mem[288 ] = 5'h10;
  assign mem[289 ] = 5'h00;
  assign mem[290 ] = 5'h01;
  assign mem[291 ] = 5'h10;
  assign mem[292 ] = 5'h00;
  assign mem[293 ] = 5'h04;
  assign mem[294 ] = 5'h13;
  assign mem[295 ] = 5'h12;
  assign mem[296 ] = 5'h11;
  assign mem[297 ] = 5'h10;
  assign mem[298 ] = 5'h00;
  assign mem[299 ] = 5'h01;
  assign mem[300 ] = 5'h10;
  assign mem[301 ] = 5'h00;
  assign mem[302 ] = 5'h02;
  assign mem[303 ] = 5'h11;
  assign mem[304 ] = 5'h10;
  assign mem[305 ] = 5'h00;
  assign mem[306 ] = 5'h01;
  assign mem[307 ] = 5'h10;
  assign mem[308 ] = 5'h00;
  assign mem[309 ] = 5'h03;
  assign mem[310 ] = 5'h12;
  assign mem[311 ] = 5'h11;
  assign mem[312 ] = 5'h10;
  assign mem[313 ] = 5'h00;
  assign mem[314 ] = 5'h01;
  assign mem[315 ] = 5'h10;
  assign mem[316 ] = 5'h00;
  assign mem[317 ] = 5'h02;
  assign mem[318 ] = 5'h11;
  assign mem[319 ] = 5'h10;
  assign mem[320 ] = 5'h00;
  assign mem[321 ] = 5'h01;
  assign mem[322 ] = 5'h10;
  assign mem[323 ] = 5'h00;
  assign mem[324 ] = 5'h05;
  assign mem[325 ] = 5'h14;
  assign mem[326 ] = 5'h13;
  assign mem[327 ] = 5'h12;
  assign mem[328 ] = 5'h11;
  assign mem[329 ] = 5'h10;
  assign mem[330 ] = 5'h00;
  assign mem[331 ] = 5'h01;
  assign mem[332 ] = 5'h10;
  assign mem[333 ] = 5'h00;
  assign mem[334 ] = 5'h02;
  assign mem[335 ] = 5'h11;
  assign mem[336 ] = 5'h10;
  assign mem[337 ] = 5'h00;
  assign mem[338 ] = 5'h01;
  assign mem[339 ] = 5'h10;
  assign mem[340 ] = 5'h00;
  assign mem[341 ] = 5'h03;
  assign mem[342 ] = 5'h12;
  assign mem[343 ] = 5'h11;
  assign mem[344 ] = 5'h10;
  assign mem[345 ] = 5'h00;
  assign mem[346 ] = 5'h01;
  assign mem[347 ] = 5'h10;
  assign mem[348 ] = 5'h00;
  assign mem[349 ] = 5'h02;
  assign mem[350 ] = 5'h11;
  assign mem[351 ] = 5'h10;
  assign mem[352 ] = 5'h00;
  assign mem[353 ] = 5'h01;
  assign mem[354 ] = 5'h10;
  assign mem[355 ] = 5'h00;
  assign mem[356 ] = 5'h04;
  assign mem[357 ] = 5'h13;
  assign mem[358 ] = 5'h12;
  assign mem[359 ] = 5'h11;
  assign mem[360 ] = 5'h10;
  assign mem[361 ] = 5'h00;
  assign mem[362 ] = 5'h01;
  assign mem[363 ] = 5'h10;
  assign mem[364 ] = 5'h00;
  assign mem[365 ] = 5'h02;
  assign mem[366 ] = 5'h11;
  assign mem[367 ] = 5'h10;
  assign mem[368 ] = 5'h00;
  assign mem[369 ] = 5'h01;
  assign mem[370 ] = 5'h10;
  assign mem[371 ] = 5'h00;
  assign mem[372 ] = 5'h03;
  assign mem[373 ] = 5'h12;
  assign mem[374 ] = 5'h11;
  assign mem[375 ] = 5'h10;
  assign mem[376 ] = 5'h00;
  assign mem[377 ] = 5'h01;
  assign mem[378 ] = 5'h10;
  assign mem[379 ] = 5'h00;
  assign mem[380 ] = 5'h02;
  assign mem[381 ] = 5'h11;
  assign mem[382 ] = 5'h10;
  assign mem[383 ] = 5'h00;
  assign mem[384 ] = 5'h01;
  assign mem[385 ] = 5'h10;
  assign mem[386 ] = 5'h00;
  assign mem[387 ] = 5'h06;
  assign mem[388 ] = 5'h15;
  assign mem[389 ] = 5'h14;
  assign mem[390 ] = 5'h13;
  assign mem[391 ] = 5'h12;
  assign mem[392 ] = 5'h11;
  assign mem[393 ] = 5'h10;
  assign mem[394 ] = 5'h00;
  assign mem[395 ] = 5'h01;
  assign mem[396 ] = 5'h10;
  assign mem[397 ] = 5'h00;
  assign mem[398 ] = 5'h02;
  assign mem[399 ] = 5'h11;
  assign mem[400 ] = 5'h10;
  assign mem[401 ] = 5'h00;
  assign mem[402 ] = 5'h01;
  assign mem[403 ] = 5'h10;
  assign mem[404 ] = 5'h00;
  assign mem[405 ] = 5'h03;
  assign mem[406 ] = 5'h12;
  assign mem[407 ] = 5'h11;
  assign mem[408 ] = 5'h10;
  assign mem[409 ] = 5'h00;
  assign mem[410 ] = 5'h01;
  assign mem[411 ] = 5'h10;
  assign mem[412 ] = 5'h00;
  assign mem[413 ] = 5'h02;
  assign mem[414 ] = 5'h11;
  assign mem[415 ] = 5'h10;
  assign mem[416 ] = 5'h00;
  assign mem[417 ] = 5'h01;
  assign mem[418 ] = 5'h10;
  assign mem[419 ] = 5'h00;
  assign mem[420 ] = 5'h04;
  assign mem[421 ] = 5'h13;
  assign mem[422 ] = 5'h12;
  assign mem[423 ] = 5'h11;
  assign mem[424 ] = 5'h10;
  assign mem[425 ] = 5'h00;
  assign mem[426 ] = 5'h01;
  assign mem[427 ] = 5'h10;
  assign mem[428 ] = 5'h00;
  assign mem[429 ] = 5'h02;
  assign mem[430 ] = 5'h11;
  assign mem[431 ] = 5'h10;
  assign mem[432 ] = 5'h00;
  assign mem[433 ] = 5'h01;
  assign mem[434 ] = 5'h10;
  assign mem[435 ] = 5'h00;
  assign mem[436 ] = 5'h03;
  assign mem[437 ] = 5'h12;
  assign mem[438 ] = 5'h11;
  assign mem[439 ] = 5'h10;
  assign mem[440 ] = 5'h00;
  assign mem[441 ] = 5'h01;
  assign mem[442 ] = 5'h10;
  assign mem[443 ] = 5'h00;
  assign mem[444 ] = 5'h02;
  assign mem[445 ] = 5'h11;
  assign mem[446 ] = 5'h10;
  assign mem[447 ] = 5'h00;
  assign mem[448 ] = 5'h01;
  assign mem[449 ] = 5'h10;
  assign mem[450 ] = 5'h00;
  assign mem[451 ] = 5'h05;
  assign mem[452 ] = 5'h14;
  assign mem[453 ] = 5'h13;
  assign mem[454 ] = 5'h12;
  assign mem[455 ] = 5'h11;
  assign mem[456 ] = 5'h10;
  assign mem[457 ] = 5'h00;
  assign mem[458 ] = 5'h01;
  assign mem[459 ] = 5'h10;
  assign mem[460 ] = 5'h00;
  assign mem[461 ] = 5'h02;
  assign mem[462 ] = 5'h11;
  assign mem[463 ] = 5'h10;
  assign mem[464 ] = 5'h00;
  assign mem[465 ] = 5'h01;
  assign mem[466 ] = 5'h10;
  assign mem[467 ] = 5'h00;
  assign mem[468 ] = 5'h03;
  assign mem[469 ] = 5'h12;
  assign mem[470 ] = 5'h11;
  assign mem[471 ] = 5'h10;
  assign mem[472 ] = 5'h00;
  assign mem[473 ] = 5'h01;
  assign mem[474 ] = 5'h10;
  assign mem[475 ] = 5'h00;
  assign mem[476 ] = 5'h02;
  assign mem[477 ] = 5'h11;
  assign mem[478 ] = 5'h10;
  assign mem[479 ] = 5'h00;
  assign mem[480 ] = 5'h01;
  assign mem[481 ] = 5'h10;
  assign mem[482 ] = 5'h00;
  assign mem[483 ] = 5'h04;
  assign mem[484 ] = 5'h13;
  assign mem[485 ] = 5'h12;
  assign mem[486 ] = 5'h11;
  assign mem[487 ] = 5'h10;
  assign mem[488 ] = 5'h00;
  assign mem[489 ] = 5'h01;
  assign mem[490 ] = 5'h10;
  assign mem[491 ] = 5'h00;
  assign mem[492 ] = 5'h02;
  assign mem[493 ] = 5'h11;
  assign mem[494 ] = 5'h10;
  assign mem[495 ] = 5'h00;
  assign mem[496 ] = 5'h01;
  assign mem[497 ] = 5'h10;
  assign mem[498 ] = 5'h00;
  assign mem[499 ] = 5'h03;
  assign mem[500 ] = 5'h12;
  assign mem[501 ] = 5'h11;
  assign mem[502 ] = 5'h10;
  assign mem[503 ] = 5'h00;
  assign mem[504 ] = 5'h01;
  assign mem[505 ] = 5'h10;
  assign mem[506 ] = 5'h00;
  assign mem[507 ] = 5'h02;
  assign mem[508 ] = 5'h11;
  assign mem[509 ] = 5'h10;
  assign mem[510 ] = 5'h00;
  assign mem[511 ] = 5'h01;
  assign mem[512 ] = 5'h10;
  assign mem[513 ] = 5'h00;
  assign mem[514 ] = 5'h08;
  assign mem[515 ] = 5'h17;
  assign mem[516 ] = 5'h16;
  assign mem[517 ] = 5'h15;
  assign mem[518 ] = 5'h14;
  assign mem[519 ] = 5'h13;
  assign mem[520 ] = 5'h12;
  assign mem[521 ] = 5'h11;
  assign mem[522 ] = 5'h10;
  assign mem[523 ] = 5'h00;
  assign mem[524 ] = 5'h01;
  assign mem[525 ] = 5'h10;
  assign mem[526 ] = 5'h00;
  assign mem[527 ] = 5'h02;
  assign mem[528 ] = 5'h11;
  assign mem[529 ] = 5'h10;
  assign mem[530 ] = 5'h00;
  assign mem[531 ] = 5'h01;
  assign mem[532 ] = 5'h10;
  assign mem[533 ] = 5'h00;
  assign mem[534 ] = 5'h03;
  assign mem[535 ] = 5'h12;
  assign mem[536 ] = 5'h11;
  assign mem[537 ] = 5'h10;
  assign mem[538 ] = 5'h00;
  assign mem[539 ] = 5'h01;
  assign mem[540 ] = 5'h10;
  assign mem[541 ] = 5'h00;
  assign mem[542 ] = 5'h02;
  assign mem[543 ] = 5'h11;
  assign mem[544 ] = 5'h10;
  assign mem[545 ] = 5'h00;
  assign mem[546 ] = 5'h01;
  assign mem[547 ] = 5'h10;
  assign mem[548 ] = 5'h00;
  assign mem[549 ] = 5'h04;
  assign mem[550 ] = 5'h13;
  assign mem[551 ] = 5'h12;
  assign mem[552 ] = 5'h11;
  assign mem[553 ] = 5'h10;
  assign mem[554 ] = 5'h00;
  assign mem[555 ] = 5'h01;
  assign mem[556 ] = 5'h10;
  assign mem[557 ] = 5'h00;
  assign mem[558 ] = 5'h02;
  assign mem[559 ] = 5'h11;
  assign mem[560 ] = 5'h10;
  assign mem[561 ] = 5'h00;
  assign mem[562 ] = 5'h01;
  assign mem[563 ] = 5'h10;
  assign mem[564 ] = 5'h00;
  assign mem[565 ] = 5'h03;
  assign mem[566 ] = 5'h12;
  assign mem[567 ] = 5'h11;
  assign mem[568 ] = 5'h10;
  assign mem[569 ] = 5'h00;
  assign mem[570 ] = 5'h01;
  assign mem[571 ] = 5'h10;
  assign mem[572 ] = 5'h00;
  assign mem[573 ] = 5'h02;
  assign mem[574 ] = 5'h11;
  assign mem[575 ] = 5'h10;
  assign mem[576 ] = 5'h00;
  assign mem[577 ] = 5'h01;
  assign mem[578 ] = 5'h10;
  assign mem[579 ] = 5'h00;
  assign mem[580 ] = 5'h05;
  assign mem[581 ] = 5'h14;
  assign mem[582 ] = 5'h13;
  assign mem[583 ] = 5'h12;
  assign mem[584 ] = 5'h11;
  assign mem[585 ] = 5'h10;
  assign mem[586 ] = 5'h00;
  assign mem[587 ] = 5'h01;
  assign mem[588 ] = 5'h10;
  assign mem[589 ] = 5'h00;
  assign mem[590 ] = 5'h02;
  assign mem[591 ] = 5'h11;
  assign mem[592 ] = 5'h10;
  assign mem[593 ] = 5'h00;
  assign mem[594 ] = 5'h01;
  assign mem[595 ] = 5'h10;
  assign mem[596 ] = 5'h00;
  assign mem[597 ] = 5'h03;
  assign mem[598 ] = 5'h12;
  assign mem[599 ] = 5'h11;
  assign mem[600 ] = 5'h10;
  assign mem[601 ] = 5'h00;
  assign mem[602 ] = 5'h01;
  assign mem[603 ] = 5'h10;
  assign mem[604 ] = 5'h00;
  assign mem[605 ] = 5'h02;
  assign mem[606 ] = 5'h11;
  assign mem[607 ] = 5'h10;
  assign mem[608 ] = 5'h00;
  assign mem[609 ] = 5'h01;
  assign mem[610 ] = 5'h10;
  assign mem[611 ] = 5'h00;
  assign mem[612 ] = 5'h04;
  assign mem[613 ] = 5'h13;
  assign mem[614 ] = 5'h12;
  assign mem[615 ] = 5'h11;
  assign mem[616 ] = 5'h10;
  assign mem[617 ] = 5'h00;
  assign mem[618 ] = 5'h01;
  assign mem[619 ] = 5'h10;
  assign mem[620 ] = 5'h00;
  assign mem[621 ] = 5'h02;
  assign mem[622 ] = 5'h11;
  assign mem[623 ] = 5'h10;
  assign mem[624 ] = 5'h00;
  assign mem[625 ] = 5'h01;
  assign mem[626 ] = 5'h10;
  assign mem[627 ] = 5'h00;
  assign mem[628 ] = 5'h03;
  assign mem[629 ] = 5'h12;
  assign mem[630 ] = 5'h11;
  assign mem[631 ] = 5'h10;
  assign mem[632 ] = 5'h00;
  assign mem[633 ] = 5'h01;
  assign mem[634 ] = 5'h10;
  assign mem[635 ] = 5'h00;
  assign mem[636 ] = 5'h02;
  assign mem[637 ] = 5'h11;
  assign mem[638 ] = 5'h10;
  assign mem[639 ] = 5'h00;
  assign mem[640 ] = 5'h01;
  assign mem[641 ] = 5'h10;
  assign mem[642 ] = 5'h00;
  assign mem[643 ] = 5'h06;
  assign mem[644 ] = 5'h15;
  assign mem[645 ] = 5'h14;
  assign mem[646 ] = 5'h13;
  assign mem[647 ] = 5'h12;
  assign mem[648 ] = 5'h11;
  assign mem[649 ] = 5'h10;
  assign mem[650 ] = 5'h00;
  assign mem[651 ] = 5'h01;
  assign mem[652 ] = 5'h10;
  assign mem[653 ] = 5'h00;
  assign mem[654 ] = 5'h02;
  assign mem[655 ] = 5'h11;
  assign mem[656 ] = 5'h10;
  assign mem[657 ] = 5'h00;
  assign mem[658 ] = 5'h01;
  assign mem[659 ] = 5'h10;
  assign mem[660 ] = 5'h00;
  assign mem[661 ] = 5'h03;
  assign mem[662 ] = 5'h12;
  assign mem[663 ] = 5'h11;
  assign mem[664 ] = 5'h10;
  assign mem[665 ] = 5'h00;
  assign mem[666 ] = 5'h01;
  assign mem[667 ] = 5'h10;
  assign mem[668 ] = 5'h00;
  assign mem[669 ] = 5'h02;
  assign mem[670 ] = 5'h11;
  assign mem[671 ] = 5'h10;
  assign mem[672 ] = 5'h00;
  assign mem[673 ] = 5'h01;
  assign mem[674 ] = 5'h10;
  assign mem[675 ] = 5'h00;
  assign mem[676 ] = 5'h04;
  assign mem[677 ] = 5'h13;
  assign mem[678 ] = 5'h12;
  assign mem[679 ] = 5'h11;
  assign mem[680 ] = 5'h10;
  assign mem[681 ] = 5'h00;
  assign mem[682 ] = 5'h01;
  assign mem[683 ] = 5'h10;
  assign mem[684 ] = 5'h00;
  assign mem[685 ] = 5'h02;
  assign mem[686 ] = 5'h11;
  assign mem[687 ] = 5'h10;
  assign mem[688 ] = 5'h00;
  assign mem[689 ] = 5'h01;
  assign mem[690 ] = 5'h10;
  assign mem[691 ] = 5'h00;
  assign mem[692 ] = 5'h03;
  assign mem[693 ] = 5'h12;
  assign mem[694 ] = 5'h11;
  assign mem[695 ] = 5'h10;
  assign mem[696 ] = 5'h00;
  assign mem[697 ] = 5'h01;
  assign mem[698 ] = 5'h10;
  assign mem[699 ] = 5'h00;
  assign mem[700 ] = 5'h02;
  assign mem[701 ] = 5'h11;
  assign mem[702 ] = 5'h10;
  assign mem[703 ] = 5'h00;
  assign mem[704 ] = 5'h01;
  assign mem[705 ] = 5'h10;
  assign mem[706 ] = 5'h00;
  assign mem[707 ] = 5'h05;
  assign mem[708 ] = 5'h14;
  assign mem[709 ] = 5'h13;
  assign mem[710 ] = 5'h12;
  assign mem[711 ] = 5'h11;
  assign mem[712 ] = 5'h10;
  assign mem[713 ] = 5'h00;
  assign mem[714 ] = 5'h01;
  assign mem[715 ] = 5'h10;
  assign mem[716 ] = 5'h00;
  assign mem[717 ] = 5'h02;
  assign mem[718 ] = 5'h11;
  assign mem[719 ] = 5'h10;
  assign mem[720 ] = 5'h00;
  assign mem[721 ] = 5'h01;
  assign mem[722 ] = 5'h10;
  assign mem[723 ] = 5'h00;
  assign mem[724 ] = 5'h03;
  assign mem[725 ] = 5'h12;
  assign mem[726 ] = 5'h11;
  assign mem[727 ] = 5'h10;
  assign mem[728 ] = 5'h00;
  assign mem[729 ] = 5'h01;
  assign mem[730 ] = 5'h10;
  assign mem[731 ] = 5'h00;
  assign mem[732 ] = 5'h02;
  assign mem[733 ] = 5'h11;
  assign mem[734 ] = 5'h10;
  assign mem[735 ] = 5'h00;
  assign mem[736 ] = 5'h01;
  assign mem[737 ] = 5'h10;
  assign mem[738 ] = 5'h00;
  assign mem[739 ] = 5'h04;
  assign mem[740 ] = 5'h13;
  assign mem[741 ] = 5'h12;
  assign mem[742 ] = 5'h11;
  assign mem[743 ] = 5'h10;
  assign mem[744 ] = 5'h00;
  assign mem[745 ] = 5'h01;
  assign mem[746 ] = 5'h10;
  assign mem[747 ] = 5'h00;
  assign mem[748 ] = 5'h02;
  assign mem[749 ] = 5'h11;
  assign mem[750 ] = 5'h10;
  assign mem[751 ] = 5'h00;
  assign mem[752 ] = 5'h01;
  assign mem[753 ] = 5'h10;
  assign mem[754 ] = 5'h00;
  assign mem[755 ] = 5'h03;
  assign mem[756 ] = 5'h12;
  assign mem[757 ] = 5'h11;
  assign mem[758 ] = 5'h10;
  assign mem[759 ] = 5'h00;
  assign mem[760 ] = 5'h01;
  assign mem[761 ] = 5'h10;
  assign mem[762 ] = 5'h00;
  assign mem[763 ] = 5'h02;
  assign mem[764 ] = 5'h11;
  assign mem[765 ] = 5'h10;
  assign mem[766 ] = 5'h00;
  assign mem[767 ] = 5'h01;
  assign mem[768 ] = 5'h10;
  assign mem[769 ] = 5'h00;
  assign mem[770 ] = 5'h07;
  assign mem[771 ] = 5'h16;
  assign mem[772 ] = 5'h15;
  assign mem[773 ] = 5'h14;
  assign mem[774 ] = 5'h13;
  assign mem[775 ] = 5'h12;
  assign mem[776 ] = 5'h11;
  assign mem[777 ] = 5'h10;
  assign mem[778 ] = 5'h00;
  assign mem[779 ] = 5'h01;
  assign mem[780 ] = 5'h10;
  assign mem[781 ] = 5'h00;
  assign mem[782 ] = 5'h02;
  assign mem[783 ] = 5'h11;
  assign mem[784 ] = 5'h10;
  assign mem[785 ] = 5'h00;
  assign mem[786 ] = 5'h01;
  assign mem[787 ] = 5'h10;
  assign mem[788 ] = 5'h00;
  assign mem[789 ] = 5'h03;
  assign mem[790 ] = 5'h12;
  assign mem[791 ] = 5'h11;
  assign mem[792 ] = 5'h10;
  assign mem[793 ] = 5'h00;
  assign mem[794 ] = 5'h01;
  assign mem[795 ] = 5'h10;
  assign mem[796 ] = 5'h00;
  assign mem[797 ] = 5'h02;
  assign mem[798 ] = 5'h11;
  assign mem[799 ] = 5'h10;
  assign mem[800 ] = 5'h00;
  assign mem[801 ] = 5'h01;
  assign mem[802 ] = 5'h10;
  assign mem[803 ] = 5'h00;
  assign mem[804 ] = 5'h04;
  assign mem[805 ] = 5'h13;
  assign mem[806 ] = 5'h12;
  assign mem[807 ] = 5'h11;
  assign mem[808 ] = 5'h10;
  assign mem[809 ] = 5'h00;
  assign mem[810 ] = 5'h01;
  assign mem[811 ] = 5'h10;
  assign mem[812 ] = 5'h00;
  assign mem[813 ] = 5'h02;
  assign mem[814 ] = 5'h11;
  assign mem[815 ] = 5'h10;
  assign mem[816 ] = 5'h00;
  assign mem[817 ] = 5'h01;
  assign mem[818 ] = 5'h10;
  assign mem[819 ] = 5'h00;
  assign mem[820 ] = 5'h03;
  assign mem[821 ] = 5'h12;
  assign mem[822 ] = 5'h11;
  assign mem[823 ] = 5'h10;
  assign mem[824 ] = 5'h00;
  assign mem[825 ] = 5'h01;
  assign mem[826 ] = 5'h10;
  assign mem[827 ] = 5'h00;
  assign mem[828 ] = 5'h02;
  assign mem[829 ] = 5'h11;
  assign mem[830 ] = 5'h10;
  assign mem[831 ] = 5'h00;
  assign mem[832 ] = 5'h01;
  assign mem[833 ] = 5'h10;
  assign mem[834 ] = 5'h00;
  assign mem[835 ] = 5'h05;
  assign mem[836 ] = 5'h14;
  assign mem[837 ] = 5'h13;
  assign mem[838 ] = 5'h12;
  assign mem[839 ] = 5'h11;
  assign mem[840 ] = 5'h10;
  assign mem[841 ] = 5'h00;
  assign mem[842 ] = 5'h01;
  assign mem[843 ] = 5'h10;
  assign mem[844 ] = 5'h00;
  assign mem[845 ] = 5'h02;
  assign mem[846 ] = 5'h11;
  assign mem[847 ] = 5'h10;
  assign mem[848 ] = 5'h00;
  assign mem[849 ] = 5'h01;
  assign mem[850 ] = 5'h10;
  assign mem[851 ] = 5'h00;
  assign mem[852 ] = 5'h03;
  assign mem[853 ] = 5'h12;
  assign mem[854 ] = 5'h11;
  assign mem[855 ] = 5'h10;
  assign mem[856 ] = 5'h00;
  assign mem[857 ] = 5'h01;
  assign mem[858 ] = 5'h10;
  assign mem[859 ] = 5'h00;
  assign mem[860 ] = 5'h02;
  assign mem[861 ] = 5'h11;
  assign mem[862 ] = 5'h10;
  assign mem[863 ] = 5'h00;
  assign mem[864 ] = 5'h01;
  assign mem[865 ] = 5'h10;
  assign mem[866 ] = 5'h00;
  assign mem[867 ] = 5'h04;
  assign mem[868 ] = 5'h13;
  assign mem[869 ] = 5'h12;
  assign mem[870 ] = 5'h11;
  assign mem[871 ] = 5'h10;
  assign mem[872 ] = 5'h00;
  assign mem[873 ] = 5'h01;
  assign mem[874 ] = 5'h10;
  assign mem[875 ] = 5'h00;
  assign mem[876 ] = 5'h02;
  assign mem[877 ] = 5'h11;
  assign mem[878 ] = 5'h10;
  assign mem[879 ] = 5'h00;
  assign mem[880 ] = 5'h01;
  assign mem[881 ] = 5'h10;
  assign mem[882 ] = 5'h00;
  assign mem[883 ] = 5'h03;
  assign mem[884 ] = 5'h12;
  assign mem[885 ] = 5'h11;
  assign mem[886 ] = 5'h10;
  assign mem[887 ] = 5'h00;
  assign mem[888 ] = 5'h01;
  assign mem[889 ] = 5'h10;
  assign mem[890 ] = 5'h00;
  assign mem[891 ] = 5'h02;
  assign mem[892 ] = 5'h11;
  assign mem[893 ] = 5'h10;
  assign mem[894 ] = 5'h00;
  assign mem[895 ] = 5'h01;
  assign mem[896 ] = 5'h10;
  assign mem[897 ] = 5'h00;
  assign mem[898 ] = 5'h06;
  assign mem[899 ] = 5'h15;
  assign mem[900 ] = 5'h14;
  assign mem[901 ] = 5'h13;
  assign mem[902 ] = 5'h12;
  assign mem[903 ] = 5'h11;
  assign mem[904 ] = 5'h10;
  assign mem[905 ] = 5'h00;
  assign mem[906 ] = 5'h01;
  assign mem[907 ] = 5'h10;
  assign mem[908 ] = 5'h00;
  assign mem[909 ] = 5'h02;
  assign mem[910 ] = 5'h11;
  assign mem[911 ] = 5'h10;
  assign mem[912 ] = 5'h00;
  assign mem[913 ] = 5'h01;
  assign mem[914 ] = 5'h10;
  assign mem[915 ] = 5'h00;
  assign mem[916 ] = 5'h03;
  assign mem[917 ] = 5'h12;
  assign mem[918 ] = 5'h11;
  assign mem[919 ] = 5'h10;
  assign mem[920 ] = 5'h00;
  assign mem[921 ] = 5'h01;
  assign mem[922 ] = 5'h10;
  assign mem[923 ] = 5'h00;
  assign mem[924 ] = 5'h02;
  assign mem[925 ] = 5'h11;
  assign mem[926 ] = 5'h10;
  assign mem[927 ] = 5'h00;
  assign mem[928 ] = 5'h01;
  assign mem[929 ] = 5'h10;
  assign mem[930 ] = 5'h00;
  assign mem[931 ] = 5'h04;
  assign mem[932 ] = 5'h13;
  assign mem[933 ] = 5'h12;
  assign mem[934 ] = 5'h11;
  assign mem[935 ] = 5'h10;
  assign mem[936 ] = 5'h00;
  assign mem[937 ] = 5'h01;
  assign mem[938 ] = 5'h10;
  assign mem[939 ] = 5'h00;
  assign mem[940 ] = 5'h02;
  assign mem[941 ] = 5'h11;
  assign mem[942 ] = 5'h10;
  assign mem[943 ] = 5'h00;
  assign mem[944 ] = 5'h01;
  assign mem[945 ] = 5'h10;
  assign mem[946 ] = 5'h00;
  assign mem[947 ] = 5'h03;
  assign mem[948 ] = 5'h12;
  assign mem[949 ] = 5'h11;
  assign mem[950 ] = 5'h10;
  assign mem[951 ] = 5'h00;
  assign mem[952 ] = 5'h01;
  assign mem[953 ] = 5'h10;
  assign mem[954 ] = 5'h00;
  assign mem[955 ] = 5'h02;
  assign mem[956 ] = 5'h11;
  assign mem[957 ] = 5'h10;
  assign mem[958 ] = 5'h00;
  assign mem[959 ] = 5'h01;
  assign mem[960 ] = 5'h10;
  assign mem[961 ] = 5'h00;
  assign mem[962 ] = 5'h05;
  assign mem[963 ] = 5'h14;
  assign mem[964 ] = 5'h13;
  assign mem[965 ] = 5'h12;
  assign mem[966 ] = 5'h11;
  assign mem[967 ] = 5'h10;
  assign mem[968 ] = 5'h00;
  assign mem[969 ] = 5'h01;
  assign mem[970 ] = 5'h10;
  assign mem[971 ] = 5'h00;
  assign mem[972 ] = 5'h02;
  assign mem[973 ] = 5'h11;
  assign mem[974 ] = 5'h10;
  assign mem[975 ] = 5'h00;
  assign mem[976 ] = 5'h01;
  assign mem[977 ] = 5'h10;
  assign mem[978 ] = 5'h00;
  assign mem[979 ] = 5'h03;
  assign mem[980 ] = 5'h12;
  assign mem[981 ] = 5'h11;
  assign mem[982 ] = 5'h10;
  assign mem[983 ] = 5'h00;
  assign mem[984 ] = 5'h01;
  assign mem[985 ] = 5'h10;
  assign mem[986 ] = 5'h00;
  assign mem[987 ] = 5'h02;
  assign mem[988 ] = 5'h11;
  assign mem[989 ] = 5'h10;
  assign mem[990 ] = 5'h00;
  assign mem[991 ] = 5'h01;
  assign mem[992 ] = 5'h10;
  assign mem[993 ] = 5'h00;
  assign mem[994 ] = 5'h04;
  assign mem[995 ] = 5'h13;
  assign mem[996 ] = 5'h12;
  assign mem[997 ] = 5'h11;
  assign mem[998 ] = 5'h10;
  assign mem[999 ] = 5'h00;
  assign mem[1000] = 5'h01;
  assign mem[1001] = 5'h10;
  assign mem[1002] = 5'h00;
  assign mem[1003] = 5'h02;
  assign mem[1004] = 5'h11;
  assign mem[1005] = 5'h10;
  assign mem[1006] = 5'h00;
  assign mem[1007] = 5'h01;
  assign mem[1008] = 5'h10;
  assign mem[1009] = 5'h00;
  assign mem[1010] = 5'h03;
  assign mem[1011] = 5'h12;
  assign mem[1012] = 5'h11;
  assign mem[1013] = 5'h10;
  assign mem[1014] = 5'h00;
  assign mem[1015] = 5'h01;
  assign mem[1016] = 5'h10;
  assign mem[1017] = 5'h00;
  assign mem[1018] = 5'h02;
  assign mem[1019] = 5'h11;
  assign mem[1020] = 5'h10;
  assign mem[1021] = 5'h00;
  assign mem[1022] = 5'h01;
  assign mem[1023] = 5'h10;
  assign mem[1024] = 5'h00;
  assign mem[1025] = 5'h09;
  assign mem[1026] = 5'h18;
  assign mem[1027] = 5'h17;
  assign mem[1028] = 5'h16;
  assign mem[1029] = 5'h15;
  assign mem[1030] = 5'h14;
  assign mem[1031] = 5'h13;
  assign mem[1032] = 5'h12;
  assign mem[1033] = 5'h11;
  assign mem[1034] = 5'h10;
  assign mem[1035] = 5'h00;
  assign mem[1036] = 5'h01;
  assign mem[1037] = 5'h10;
  assign mem[1038] = 5'h00;
  assign mem[1039] = 5'h02;
  assign mem[1040] = 5'h11;
  assign mem[1041] = 5'h10;
  assign mem[1042] = 5'h00;
  assign mem[1043] = 5'h01;
  assign mem[1044] = 5'h10;
  assign mem[1045] = 5'h00;
  assign mem[1046] = 5'h03;
  assign mem[1047] = 5'h12;
  assign mem[1048] = 5'h11;
  assign mem[1049] = 5'h10;
  assign mem[1050] = 5'h00;
  assign mem[1051] = 5'h01;
  assign mem[1052] = 5'h10;
  assign mem[1053] = 5'h00;
  assign mem[1054] = 5'h02;
  assign mem[1055] = 5'h11;
  assign mem[1056] = 5'h10;
  assign mem[1057] = 5'h00;
  assign mem[1058] = 5'h01;
  assign mem[1059] = 5'h10;
  assign mem[1060] = 5'h00;
  assign mem[1061] = 5'h04;
  assign mem[1062] = 5'h13;
  assign mem[1063] = 5'h12;
  assign mem[1064] = 5'h11;
  assign mem[1065] = 5'h10;
  assign mem[1066] = 5'h00;
  assign mem[1067] = 5'h01;
  assign mem[1068] = 5'h10;
  assign mem[1069] = 5'h00;
  assign mem[1070] = 5'h02;
  assign mem[1071] = 5'h11;
  assign mem[1072] = 5'h10;
  assign mem[1073] = 5'h00;
  assign mem[1074] = 5'h01;
  assign mem[1075] = 5'h10;
  assign mem[1076] = 5'h00;
  assign mem[1077] = 5'h03;
  assign mem[1078] = 5'h12;
  assign mem[1079] = 5'h11;
  assign mem[1080] = 5'h10;
  assign mem[1081] = 5'h00;
  assign mem[1082] = 5'h01;
  assign mem[1083] = 5'h10;
  assign mem[1084] = 5'h00;
  assign mem[1085] = 5'h02;
  assign mem[1086] = 5'h11;
  assign mem[1087] = 5'h10;
  assign mem[1088] = 5'h00;
  assign mem[1089] = 5'h01;
  assign mem[1090] = 5'h10;
  assign mem[1091] = 5'h00;
  assign mem[1092] = 5'h05;
  assign mem[1093] = 5'h14;
  assign mem[1094] = 5'h13;
  assign mem[1095] = 5'h12;
  assign mem[1096] = 5'h11;
  assign mem[1097] = 5'h10;
  assign mem[1098] = 5'h00;
  assign mem[1099] = 5'h01;
  assign mem[1100] = 5'h10;
  assign mem[1101] = 5'h00;
  assign mem[1102] = 5'h02;
  assign mem[1103] = 5'h11;
  assign mem[1104] = 5'h10;
  assign mem[1105] = 5'h00;
  assign mem[1106] = 5'h01;
  assign mem[1107] = 5'h10;
  assign mem[1108] = 5'h00;
  assign mem[1109] = 5'h03;
  assign mem[1110] = 5'h12;
  assign mem[1111] = 5'h11;
  assign mem[1112] = 5'h10;
  assign mem[1113] = 5'h00;
  assign mem[1114] = 5'h01;
  assign mem[1115] = 5'h10;
  assign mem[1116] = 5'h00;
  assign mem[1117] = 5'h02;
  assign mem[1118] = 5'h11;
  assign mem[1119] = 5'h10;
  assign mem[1120] = 5'h00;
  assign mem[1121] = 5'h01;
  assign mem[1122] = 5'h10;
  assign mem[1123] = 5'h00;
  assign mem[1124] = 5'h04;
  assign mem[1125] = 5'h13;
  assign mem[1126] = 5'h12;
  assign mem[1127] = 5'h11;
  assign mem[1128] = 5'h10;
  assign mem[1129] = 5'h00;
  assign mem[1130] = 5'h01;
  assign mem[1131] = 5'h10;
  assign mem[1132] = 5'h00;
  assign mem[1133] = 5'h02;
  assign mem[1134] = 5'h11;
  assign mem[1135] = 5'h10;
  assign mem[1136] = 5'h00;
  assign mem[1137] = 5'h01;
  assign mem[1138] = 5'h10;
  assign mem[1139] = 5'h00;
  assign mem[1140] = 5'h03;
  assign mem[1141] = 5'h12;
  assign mem[1142] = 5'h11;
  assign mem[1143] = 5'h10;
  assign mem[1144] = 5'h00;
  assign mem[1145] = 5'h01;
  assign mem[1146] = 5'h10;
  assign mem[1147] = 5'h00;
  assign mem[1148] = 5'h02;
  assign mem[1149] = 5'h11;
  assign mem[1150] = 5'h10;
  assign mem[1151] = 5'h00;
  assign mem[1152] = 5'h01;
  assign mem[1153] = 5'h10;
  assign mem[1154] = 5'h00;
  assign mem[1155] = 5'h06;
  assign mem[1156] = 5'h15;
  assign mem[1157] = 5'h14;
  assign mem[1158] = 5'h13;
  assign mem[1159] = 5'h12;
  assign mem[1160] = 5'h11;
  assign mem[1161] = 5'h10;
  assign mem[1162] = 5'h00;
  assign mem[1163] = 5'h01;
  assign mem[1164] = 5'h10;
  assign mem[1165] = 5'h00;
  assign mem[1166] = 5'h02;
  assign mem[1167] = 5'h11;
  assign mem[1168] = 5'h10;
  assign mem[1169] = 5'h00;
  assign mem[1170] = 5'h01;
  assign mem[1171] = 5'h10;
  assign mem[1172] = 5'h00;
  assign mem[1173] = 5'h03;
  assign mem[1174] = 5'h12;
  assign mem[1175] = 5'h11;
  assign mem[1176] = 5'h10;
  assign mem[1177] = 5'h00;
  assign mem[1178] = 5'h01;
  assign mem[1179] = 5'h10;
  assign mem[1180] = 5'h00;
  assign mem[1181] = 5'h02;
  assign mem[1182] = 5'h11;
  assign mem[1183] = 5'h10;
  assign mem[1184] = 5'h00;
  assign mem[1185] = 5'h01;
  assign mem[1186] = 5'h10;
  assign mem[1187] = 5'h00;
  assign mem[1188] = 5'h04;
  assign mem[1189] = 5'h13;
  assign mem[1190] = 5'h12;
  assign mem[1191] = 5'h11;
  assign mem[1192] = 5'h10;
  assign mem[1193] = 5'h00;
  assign mem[1194] = 5'h01;
  assign mem[1195] = 5'h10;
  assign mem[1196] = 5'h00;
  assign mem[1197] = 5'h02;
  assign mem[1198] = 5'h11;
  assign mem[1199] = 5'h10;
  assign mem[1200] = 5'h00;
  assign mem[1201] = 5'h01;
  assign mem[1202] = 5'h10;
  assign mem[1203] = 5'h00;
  assign mem[1204] = 5'h03;
  assign mem[1205] = 5'h12;
  assign mem[1206] = 5'h11;
  assign mem[1207] = 5'h10;
  assign mem[1208] = 5'h00;
  assign mem[1209] = 5'h01;
  assign mem[1210] = 5'h10;
  assign mem[1211] = 5'h00;
  assign mem[1212] = 5'h02;
  assign mem[1213] = 5'h11;
  assign mem[1214] = 5'h10;
  assign mem[1215] = 5'h00;
  assign mem[1216] = 5'h01;
  assign mem[1217] = 5'h10;
  assign mem[1218] = 5'h00;
  assign mem[1219] = 5'h05;
  assign mem[1220] = 5'h14;
  assign mem[1221] = 5'h13;
  assign mem[1222] = 5'h12;
  assign mem[1223] = 5'h11;
  assign mem[1224] = 5'h10;
  assign mem[1225] = 5'h00;
  assign mem[1226] = 5'h01;
  assign mem[1227] = 5'h10;
  assign mem[1228] = 5'h00;
  assign mem[1229] = 5'h02;
  assign mem[1230] = 5'h11;
  assign mem[1231] = 5'h10;
  assign mem[1232] = 5'h00;
  assign mem[1233] = 5'h01;
  assign mem[1234] = 5'h10;
  assign mem[1235] = 5'h00;
  assign mem[1236] = 5'h03;
  assign mem[1237] = 5'h12;
  assign mem[1238] = 5'h11;
  assign mem[1239] = 5'h10;
  assign mem[1240] = 5'h00;
  assign mem[1241] = 5'h01;
  assign mem[1242] = 5'h10;
  assign mem[1243] = 5'h00;
  assign mem[1244] = 5'h02;
  assign mem[1245] = 5'h11;
  assign mem[1246] = 5'h10;
  assign mem[1247] = 5'h00;
  assign mem[1248] = 5'h01;
  assign mem[1249] = 5'h10;
  assign mem[1250] = 5'h00;
  assign mem[1251] = 5'h04;
  assign mem[1252] = 5'h13;
  assign mem[1253] = 5'h12;
  assign mem[1254] = 5'h11;
  assign mem[1255] = 5'h10;
  assign mem[1256] = 5'h00;
  assign mem[1257] = 5'h01;
  assign mem[1258] = 5'h10;
  assign mem[1259] = 5'h00;
  assign mem[1260] = 5'h02;
  assign mem[1261] = 5'h11;
  assign mem[1262] = 5'h10;
  assign mem[1263] = 5'h00;
  assign mem[1264] = 5'h01;
  assign mem[1265] = 5'h10;
  assign mem[1266] = 5'h00;
  assign mem[1267] = 5'h03;
  assign mem[1268] = 5'h12;
  assign mem[1269] = 5'h11;
  assign mem[1270] = 5'h10;
  assign mem[1271] = 5'h00;
  assign mem[1272] = 5'h01;
  assign mem[1273] = 5'h10;
  assign mem[1274] = 5'h00;
  assign mem[1275] = 5'h02;
  assign mem[1276] = 5'h11;
  assign mem[1277] = 5'h10;
  assign mem[1278] = 5'h00;
  assign mem[1279] = 5'h01;
  assign mem[1280] = 5'h10;
  assign mem[1281] = 5'h00;
  assign mem[1282] = 5'h07;
  assign mem[1283] = 5'h16;
  assign mem[1284] = 5'h15;
  assign mem[1285] = 5'h14;
  assign mem[1286] = 5'h13;
  assign mem[1287] = 5'h12;
  assign mem[1288] = 5'h11;
  assign mem[1289] = 5'h10;
  assign mem[1290] = 5'h00;
  assign mem[1291] = 5'h01;
  assign mem[1292] = 5'h10;
  assign mem[1293] = 5'h00;
  assign mem[1294] = 5'h02;
  assign mem[1295] = 5'h11;
  assign mem[1296] = 5'h10;
  assign mem[1297] = 5'h00;
  assign mem[1298] = 5'h01;
  assign mem[1299] = 5'h10;
  assign mem[1300] = 5'h00;
  assign mem[1301] = 5'h03;
  assign mem[1302] = 5'h12;
  assign mem[1303] = 5'h11;
  assign mem[1304] = 5'h10;
  assign mem[1305] = 5'h00;
  assign mem[1306] = 5'h01;
  assign mem[1307] = 5'h10;
  assign mem[1308] = 5'h00;
  assign mem[1309] = 5'h02;
  assign mem[1310] = 5'h11;
  assign mem[1311] = 5'h10;
  assign mem[1312] = 5'h00;
  assign mem[1313] = 5'h01;
  assign mem[1314] = 5'h10;
  assign mem[1315] = 5'h00;
  assign mem[1316] = 5'h04;
  assign mem[1317] = 5'h13;
  assign mem[1318] = 5'h12;
  assign mem[1319] = 5'h11;
  assign mem[1320] = 5'h10;
  assign mem[1321] = 5'h00;
  assign mem[1322] = 5'h01;
  assign mem[1323] = 5'h10;
  assign mem[1324] = 5'h00;
  assign mem[1325] = 5'h02;
  assign mem[1326] = 5'h11;
  assign mem[1327] = 5'h10;
  assign mem[1328] = 5'h00;
  assign mem[1329] = 5'h01;
  assign mem[1330] = 5'h10;
  assign mem[1331] = 5'h00;
  assign mem[1332] = 5'h03;
  assign mem[1333] = 5'h12;
  assign mem[1334] = 5'h11;
  assign mem[1335] = 5'h10;
  assign mem[1336] = 5'h00;
  assign mem[1337] = 5'h01;
  assign mem[1338] = 5'h10;
  assign mem[1339] = 5'h00;
  assign mem[1340] = 5'h02;
  assign mem[1341] = 5'h11;
  assign mem[1342] = 5'h10;
  assign mem[1343] = 5'h00;
  assign mem[1344] = 5'h01;
  assign mem[1345] = 5'h10;
  assign mem[1346] = 5'h00;
  assign mem[1347] = 5'h05;
  assign mem[1348] = 5'h14;
  assign mem[1349] = 5'h13;
  assign mem[1350] = 5'h12;
  assign mem[1351] = 5'h11;
  assign mem[1352] = 5'h10;
  assign mem[1353] = 5'h00;
  assign mem[1354] = 5'h01;
  assign mem[1355] = 5'h10;
  assign mem[1356] = 5'h00;
  assign mem[1357] = 5'h02;
  assign mem[1358] = 5'h11;
  assign mem[1359] = 5'h10;
  assign mem[1360] = 5'h00;
  assign mem[1361] = 5'h01;
  assign mem[1362] = 5'h10;
  assign mem[1363] = 5'h00;
  assign mem[1364] = 5'h03;
  assign mem[1365] = 5'h12;
  assign mem[1366] = 5'h11;
  assign mem[1367] = 5'h10;
  assign mem[1368] = 5'h00;
  assign mem[1369] = 5'h01;
  assign mem[1370] = 5'h10;
  assign mem[1371] = 5'h00;
  assign mem[1372] = 5'h02;
  assign mem[1373] = 5'h11;
  assign mem[1374] = 5'h10;
  assign mem[1375] = 5'h00;
  assign mem[1376] = 5'h01;
  assign mem[1377] = 5'h10;
  assign mem[1378] = 5'h00;
  assign mem[1379] = 5'h04;
  assign mem[1380] = 5'h13;
  assign mem[1381] = 5'h12;
  assign mem[1382] = 5'h11;
  assign mem[1383] = 5'h10;
  assign mem[1384] = 5'h00;
  assign mem[1385] = 5'h01;
  assign mem[1386] = 5'h10;
  assign mem[1387] = 5'h00;
  assign mem[1388] = 5'h02;
  assign mem[1389] = 5'h11;
  assign mem[1390] = 5'h10;
  assign mem[1391] = 5'h00;
  assign mem[1392] = 5'h01;
  assign mem[1393] = 5'h10;
  assign mem[1394] = 5'h00;
  assign mem[1395] = 5'h03;
  assign mem[1396] = 5'h12;
  assign mem[1397] = 5'h11;
  assign mem[1398] = 5'h10;
  assign mem[1399] = 5'h00;
  assign mem[1400] = 5'h01;
  assign mem[1401] = 5'h10;
  assign mem[1402] = 5'h00;
  assign mem[1403] = 5'h02;
  assign mem[1404] = 5'h11;
  assign mem[1405] = 5'h10;
  assign mem[1406] = 5'h00;
  assign mem[1407] = 5'h01;
  assign mem[1408] = 5'h10;
  assign mem[1409] = 5'h00;
  assign mem[1410] = 5'h06;
  assign mem[1411] = 5'h15;
  assign mem[1412] = 5'h14;
  assign mem[1413] = 5'h13;
  assign mem[1414] = 5'h12;
  assign mem[1415] = 5'h11;
  assign mem[1416] = 5'h10;
  assign mem[1417] = 5'h00;
  assign mem[1418] = 5'h01;
  assign mem[1419] = 5'h10;
  assign mem[1420] = 5'h00;
  assign mem[1421] = 5'h02;
  assign mem[1422] = 5'h11;
  assign mem[1423] = 5'h10;
  assign mem[1424] = 5'h00;
  assign mem[1425] = 5'h01;
  assign mem[1426] = 5'h10;
  assign mem[1427] = 5'h00;
  assign mem[1428] = 5'h03;
  assign mem[1429] = 5'h12;
  assign mem[1430] = 5'h11;
  assign mem[1431] = 5'h10;
  assign mem[1432] = 5'h00;
  assign mem[1433] = 5'h01;
  assign mem[1434] = 5'h10;
  assign mem[1435] = 5'h00;
  assign mem[1436] = 5'h02;
  assign mem[1437] = 5'h11;
  assign mem[1438] = 5'h10;
  assign mem[1439] = 5'h00;
  assign mem[1440] = 5'h01;
  assign mem[1441] = 5'h10;
  assign mem[1442] = 5'h00;
  assign mem[1443] = 5'h04;
  assign mem[1444] = 5'h13;
  assign mem[1445] = 5'h12;
  assign mem[1446] = 5'h11;
  assign mem[1447] = 5'h10;
  assign mem[1448] = 5'h00;
  assign mem[1449] = 5'h01;
  assign mem[1450] = 5'h10;
  assign mem[1451] = 5'h00;
  assign mem[1452] = 5'h02;
  assign mem[1453] = 5'h11;
  assign mem[1454] = 5'h10;
  assign mem[1455] = 5'h00;
  assign mem[1456] = 5'h01;
  assign mem[1457] = 5'h10;
  assign mem[1458] = 5'h00;
  assign mem[1459] = 5'h03;
  assign mem[1460] = 5'h12;
  assign mem[1461] = 5'h11;
  assign mem[1462] = 5'h10;
  assign mem[1463] = 5'h00;
  assign mem[1464] = 5'h01;
  assign mem[1465] = 5'h10;
  assign mem[1466] = 5'h00;
  assign mem[1467] = 5'h02;
  assign mem[1468] = 5'h11;
  assign mem[1469] = 5'h10;
  assign mem[1470] = 5'h00;
  assign mem[1471] = 5'h01;
  assign mem[1472] = 5'h10;
  assign mem[1473] = 5'h00;
  assign mem[1474] = 5'h05;
  assign mem[1475] = 5'h14;
  assign mem[1476] = 5'h13;
  assign mem[1477] = 5'h12;
  assign mem[1478] = 5'h11;
  assign mem[1479] = 5'h10;
  assign mem[1480] = 5'h00;
  assign mem[1481] = 5'h01;
  assign mem[1482] = 5'h10;
  assign mem[1483] = 5'h00;
  assign mem[1484] = 5'h02;
  assign mem[1485] = 5'h11;
  assign mem[1486] = 5'h10;
  assign mem[1487] = 5'h00;
  assign mem[1488] = 5'h01;
  assign mem[1489] = 5'h10;
  assign mem[1490] = 5'h00;
  assign mem[1491] = 5'h03;
  assign mem[1492] = 5'h12;
  assign mem[1493] = 5'h11;
  assign mem[1494] = 5'h10;
  assign mem[1495] = 5'h00;
  assign mem[1496] = 5'h01;
  assign mem[1497] = 5'h10;
  assign mem[1498] = 5'h00;
  assign mem[1499] = 5'h02;
  assign mem[1500] = 5'h11;
  assign mem[1501] = 5'h10;
  assign mem[1502] = 5'h00;
  assign mem[1503] = 5'h01;
  assign mem[1504] = 5'h10;
  assign mem[1505] = 5'h00;
  assign mem[1506] = 5'h04;
  assign mem[1507] = 5'h13;
  assign mem[1508] = 5'h12;
  assign mem[1509] = 5'h11;
  assign mem[1510] = 5'h10;
  assign mem[1511] = 5'h00;
  assign mem[1512] = 5'h01;
  assign mem[1513] = 5'h10;
  assign mem[1514] = 5'h00;
  assign mem[1515] = 5'h02;
  assign mem[1516] = 5'h11;
  assign mem[1517] = 5'h10;
  assign mem[1518] = 5'h00;
  assign mem[1519] = 5'h01;
  assign mem[1520] = 5'h10;
  assign mem[1521] = 5'h00;
  assign mem[1522] = 5'h03;
  assign mem[1523] = 5'h12;
  assign mem[1524] = 5'h11;
  assign mem[1525] = 5'h10;
  assign mem[1526] = 5'h00;
  assign mem[1527] = 5'h01;
  assign mem[1528] = 5'h10;
  assign mem[1529] = 5'h00;
  assign mem[1530] = 5'h02;
  assign mem[1531] = 5'h11;
  assign mem[1532] = 5'h10;
  assign mem[1533] = 5'h00;
  assign mem[1534] = 5'h01;
  assign mem[1535] = 5'h10;
  assign mem[1536] = 5'h00;
  assign mem[1537] = 5'h08;
  assign mem[1538] = 5'h17;
  assign mem[1539] = 5'h16;
  assign mem[1540] = 5'h15;
  assign mem[1541] = 5'h14;
  assign mem[1542] = 5'h13;
  assign mem[1543] = 5'h12;
  assign mem[1544] = 5'h11;
  assign mem[1545] = 5'h10;
  assign mem[1546] = 5'h00;
  assign mem[1547] = 5'h01;
  assign mem[1548] = 5'h10;
  assign mem[1549] = 5'h00;
  assign mem[1550] = 5'h02;
  assign mem[1551] = 5'h11;
  assign mem[1552] = 5'h10;
  assign mem[1553] = 5'h00;
  assign mem[1554] = 5'h01;
  assign mem[1555] = 5'h10;
  assign mem[1556] = 5'h00;
  assign mem[1557] = 5'h03;
  assign mem[1558] = 5'h12;
  assign mem[1559] = 5'h11;
  assign mem[1560] = 5'h10;
  assign mem[1561] = 5'h00;
  assign mem[1562] = 5'h01;
  assign mem[1563] = 5'h10;
  assign mem[1564] = 5'h00;
  assign mem[1565] = 5'h02;
  assign mem[1566] = 5'h11;
  assign mem[1567] = 5'h10;
  assign mem[1568] = 5'h00;
  assign mem[1569] = 5'h01;
  assign mem[1570] = 5'h10;
  assign mem[1571] = 5'h00;
  assign mem[1572] = 5'h04;
  assign mem[1573] = 5'h13;
  assign mem[1574] = 5'h12;
  assign mem[1575] = 5'h11;
  assign mem[1576] = 5'h10;
  assign mem[1577] = 5'h00;
  assign mem[1578] = 5'h01;
  assign mem[1579] = 5'h10;
  assign mem[1580] = 5'h00;
  assign mem[1581] = 5'h02;
  assign mem[1582] = 5'h11;
  assign mem[1583] = 5'h10;
  assign mem[1584] = 5'h00;
  assign mem[1585] = 5'h01;
  assign mem[1586] = 5'h10;
  assign mem[1587] = 5'h00;
  assign mem[1588] = 5'h03;
  assign mem[1589] = 5'h12;
  assign mem[1590] = 5'h11;
  assign mem[1591] = 5'h10;
  assign mem[1592] = 5'h00;
  assign mem[1593] = 5'h01;
  assign mem[1594] = 5'h10;
  assign mem[1595] = 5'h00;
  assign mem[1596] = 5'h02;
  assign mem[1597] = 5'h11;
  assign mem[1598] = 5'h10;
  assign mem[1599] = 5'h00;
  assign mem[1600] = 5'h01;
  assign mem[1601] = 5'h10;
  assign mem[1602] = 5'h00;
  assign mem[1603] = 5'h05;
  assign mem[1604] = 5'h14;
  assign mem[1605] = 5'h13;
  assign mem[1606] = 5'h12;
  assign mem[1607] = 5'h11;
  assign mem[1608] = 5'h10;
  assign mem[1609] = 5'h00;
  assign mem[1610] = 5'h01;
  assign mem[1611] = 5'h10;
  assign mem[1612] = 5'h00;
  assign mem[1613] = 5'h02;
  assign mem[1614] = 5'h11;
  assign mem[1615] = 5'h10;
  assign mem[1616] = 5'h00;
  assign mem[1617] = 5'h01;
  assign mem[1618] = 5'h10;
  assign mem[1619] = 5'h00;
  assign mem[1620] = 5'h03;
  assign mem[1621] = 5'h12;
  assign mem[1622] = 5'h11;
  assign mem[1623] = 5'h10;
  assign mem[1624] = 5'h00;
  assign mem[1625] = 5'h01;
  assign mem[1626] = 5'h10;
  assign mem[1627] = 5'h00;
  assign mem[1628] = 5'h02;
  assign mem[1629] = 5'h11;
  assign mem[1630] = 5'h10;
  assign mem[1631] = 5'h00;
  assign mem[1632] = 5'h01;
  assign mem[1633] = 5'h10;
  assign mem[1634] = 5'h00;
  assign mem[1635] = 5'h04;
  assign mem[1636] = 5'h13;
  assign mem[1637] = 5'h12;
  assign mem[1638] = 5'h11;
  assign mem[1639] = 5'h10;
  assign mem[1640] = 5'h00;
  assign mem[1641] = 5'h01;
  assign mem[1642] = 5'h10;
  assign mem[1643] = 5'h00;
  assign mem[1644] = 5'h02;
  assign mem[1645] = 5'h11;
  assign mem[1646] = 5'h10;
  assign mem[1647] = 5'h00;
  assign mem[1648] = 5'h01;
  assign mem[1649] = 5'h10;
  assign mem[1650] = 5'h00;
  assign mem[1651] = 5'h03;
  assign mem[1652] = 5'h12;
  assign mem[1653] = 5'h11;
  assign mem[1654] = 5'h10;
  assign mem[1655] = 5'h00;
  assign mem[1656] = 5'h01;
  assign mem[1657] = 5'h10;
  assign mem[1658] = 5'h00;
  assign mem[1659] = 5'h02;
  assign mem[1660] = 5'h11;
  assign mem[1661] = 5'h10;
  assign mem[1662] = 5'h00;
  assign mem[1663] = 5'h01;
  assign mem[1664] = 5'h10;
  assign mem[1665] = 5'h00;
  assign mem[1666] = 5'h06;
  assign mem[1667] = 5'h15;
  assign mem[1668] = 5'h14;
  assign mem[1669] = 5'h13;
  assign mem[1670] = 5'h12;
  assign mem[1671] = 5'h11;
  assign mem[1672] = 5'h10;
  assign mem[1673] = 5'h00;
  assign mem[1674] = 5'h01;
  assign mem[1675] = 5'h10;
  assign mem[1676] = 5'h00;
  assign mem[1677] = 5'h02;
  assign mem[1678] = 5'h11;
  assign mem[1679] = 5'h10;
  assign mem[1680] = 5'h00;
  assign mem[1681] = 5'h01;
  assign mem[1682] = 5'h10;
  assign mem[1683] = 5'h00;
  assign mem[1684] = 5'h03;
  assign mem[1685] = 5'h12;
  assign mem[1686] = 5'h11;
  assign mem[1687] = 5'h10;
  assign mem[1688] = 5'h00;
  assign mem[1689] = 5'h01;
  assign mem[1690] = 5'h10;
  assign mem[1691] = 5'h00;
  assign mem[1692] = 5'h02;
  assign mem[1693] = 5'h11;
  assign mem[1694] = 5'h10;
  assign mem[1695] = 5'h00;
  assign mem[1696] = 5'h01;
  assign mem[1697] = 5'h10;
  assign mem[1698] = 5'h00;
  assign mem[1699] = 5'h04;
  assign mem[1700] = 5'h13;
  assign mem[1701] = 5'h12;
  assign mem[1702] = 5'h11;
  assign mem[1703] = 5'h10;
  assign mem[1704] = 5'h00;
  assign mem[1705] = 5'h01;
  assign mem[1706] = 5'h10;
  assign mem[1707] = 5'h00;
  assign mem[1708] = 5'h02;
  assign mem[1709] = 5'h11;
  assign mem[1710] = 5'h10;
  assign mem[1711] = 5'h00;
  assign mem[1712] = 5'h01;
  assign mem[1713] = 5'h10;
  assign mem[1714] = 5'h00;
  assign mem[1715] = 5'h03;
  assign mem[1716] = 5'h12;
  assign mem[1717] = 5'h11;
  assign mem[1718] = 5'h10;
  assign mem[1719] = 5'h00;
  assign mem[1720] = 5'h01;
  assign mem[1721] = 5'h10;
  assign mem[1722] = 5'h00;
  assign mem[1723] = 5'h02;
  assign mem[1724] = 5'h11;
  assign mem[1725] = 5'h10;
  assign mem[1726] = 5'h00;
  assign mem[1727] = 5'h01;
  assign mem[1728] = 5'h10;
  assign mem[1729] = 5'h00;
  assign mem[1730] = 5'h05;
  assign mem[1731] = 5'h14;
  assign mem[1732] = 5'h13;
  assign mem[1733] = 5'h12;
  assign mem[1734] = 5'h11;
  assign mem[1735] = 5'h10;
  assign mem[1736] = 5'h00;
  assign mem[1737] = 5'h01;
  assign mem[1738] = 5'h10;
  assign mem[1739] = 5'h00;
  assign mem[1740] = 5'h02;
  assign mem[1741] = 5'h11;
  assign mem[1742] = 5'h10;
  assign mem[1743] = 5'h00;
  assign mem[1744] = 5'h01;
  assign mem[1745] = 5'h10;
  assign mem[1746] = 5'h00;
  assign mem[1747] = 5'h03;
  assign mem[1748] = 5'h12;
  assign mem[1749] = 5'h11;
  assign mem[1750] = 5'h10;
  assign mem[1751] = 5'h00;
  assign mem[1752] = 5'h01;
  assign mem[1753] = 5'h10;
  assign mem[1754] = 5'h00;
  assign mem[1755] = 5'h02;
  assign mem[1756] = 5'h11;
  assign mem[1757] = 5'h10;
  assign mem[1758] = 5'h00;
  assign mem[1759] = 5'h01;
  assign mem[1760] = 5'h10;
  assign mem[1761] = 5'h00;
  assign mem[1762] = 5'h04;
  assign mem[1763] = 5'h13;
  assign mem[1764] = 5'h12;
  assign mem[1765] = 5'h11;
  assign mem[1766] = 5'h10;
  assign mem[1767] = 5'h00;
  assign mem[1768] = 5'h01;
  assign mem[1769] = 5'h10;
  assign mem[1770] = 5'h00;
  assign mem[1771] = 5'h02;
  assign mem[1772] = 5'h11;
  assign mem[1773] = 5'h10;
  assign mem[1774] = 5'h00;
  assign mem[1775] = 5'h01;
  assign mem[1776] = 5'h10;
  assign mem[1777] = 5'h00;
  assign mem[1778] = 5'h03;
  assign mem[1779] = 5'h12;
  assign mem[1780] = 5'h11;
  assign mem[1781] = 5'h10;
  assign mem[1782] = 5'h00;
  assign mem[1783] = 5'h01;
  assign mem[1784] = 5'h10;
  assign mem[1785] = 5'h00;
  assign mem[1786] = 5'h02;
  assign mem[1787] = 5'h11;
  assign mem[1788] = 5'h10;
  assign mem[1789] = 5'h00;
  assign mem[1790] = 5'h01;
  assign mem[1791] = 5'h10;
  assign mem[1792] = 5'h00;
  assign mem[1793] = 5'h07;
  assign mem[1794] = 5'h16;
  assign mem[1795] = 5'h15;
  assign mem[1796] = 5'h14;
  assign mem[1797] = 5'h13;
  assign mem[1798] = 5'h12;
  assign mem[1799] = 5'h11;
  assign mem[1800] = 5'h10;
  assign mem[1801] = 5'h00;
  assign mem[1802] = 5'h01;
  assign mem[1803] = 5'h10;
  assign mem[1804] = 5'h00;
  assign mem[1805] = 5'h02;
  assign mem[1806] = 5'h11;
  assign mem[1807] = 5'h10;
  assign mem[1808] = 5'h00;
  assign mem[1809] = 5'h01;
  assign mem[1810] = 5'h10;
  assign mem[1811] = 5'h00;
  assign mem[1812] = 5'h03;
  assign mem[1813] = 5'h12;
  assign mem[1814] = 5'h11;
  assign mem[1815] = 5'h10;
  assign mem[1816] = 5'h00;
  assign mem[1817] = 5'h01;
  assign mem[1818] = 5'h10;
  assign mem[1819] = 5'h00;
  assign mem[1820] = 5'h02;
  assign mem[1821] = 5'h11;
  assign mem[1822] = 5'h10;
  assign mem[1823] = 5'h00;
  assign mem[1824] = 5'h01;
  assign mem[1825] = 5'h10;
  assign mem[1826] = 5'h00;
  assign mem[1827] = 5'h04;
  assign mem[1828] = 5'h13;
  assign mem[1829] = 5'h12;
  assign mem[1830] = 5'h11;
  assign mem[1831] = 5'h10;
  assign mem[1832] = 5'h00;
  assign mem[1833] = 5'h01;
  assign mem[1834] = 5'h10;
  assign mem[1835] = 5'h00;
  assign mem[1836] = 5'h02;
  assign mem[1837] = 5'h11;
  assign mem[1838] = 5'h10;
  assign mem[1839] = 5'h00;
  assign mem[1840] = 5'h01;
  assign mem[1841] = 5'h10;
  assign mem[1842] = 5'h00;
  assign mem[1843] = 5'h03;
  assign mem[1844] = 5'h12;
  assign mem[1845] = 5'h11;
  assign mem[1846] = 5'h10;
  assign mem[1847] = 5'h00;
  assign mem[1848] = 5'h01;
  assign mem[1849] = 5'h10;
  assign mem[1850] = 5'h00;
  assign mem[1851] = 5'h02;
  assign mem[1852] = 5'h11;
  assign mem[1853] = 5'h10;
  assign mem[1854] = 5'h00;
  assign mem[1855] = 5'h01;
  assign mem[1856] = 5'h10;
  assign mem[1857] = 5'h00;
  assign mem[1858] = 5'h05;
  assign mem[1859] = 5'h14;
  assign mem[1860] = 5'h13;
  assign mem[1861] = 5'h12;
  assign mem[1862] = 5'h11;
  assign mem[1863] = 5'h10;
  assign mem[1864] = 5'h00;
  assign mem[1865] = 5'h01;
  assign mem[1866] = 5'h10;
  assign mem[1867] = 5'h00;
  assign mem[1868] = 5'h02;
  assign mem[1869] = 5'h11;
  assign mem[1870] = 5'h10;
  assign mem[1871] = 5'h00;
  assign mem[1872] = 5'h01;
  assign mem[1873] = 5'h10;
  assign mem[1874] = 5'h00;
  assign mem[1875] = 5'h03;
  assign mem[1876] = 5'h12;
  assign mem[1877] = 5'h11;
  assign mem[1878] = 5'h10;
  assign mem[1879] = 5'h00;
  assign mem[1880] = 5'h01;
  assign mem[1881] = 5'h10;
  assign mem[1882] = 5'h00;
  assign mem[1883] = 5'h02;
  assign mem[1884] = 5'h11;
  assign mem[1885] = 5'h10;
  assign mem[1886] = 5'h00;
  assign mem[1887] = 5'h01;
  assign mem[1888] = 5'h10;
  assign mem[1889] = 5'h00;
  assign mem[1890] = 5'h04;
  assign mem[1891] = 5'h13;
  assign mem[1892] = 5'h12;
  assign mem[1893] = 5'h11;
  assign mem[1894] = 5'h10;
  assign mem[1895] = 5'h00;
  assign mem[1896] = 5'h01;
  assign mem[1897] = 5'h10;
  assign mem[1898] = 5'h00;
  assign mem[1899] = 5'h02;
  assign mem[1900] = 5'h11;
  assign mem[1901] = 5'h10;
  assign mem[1902] = 5'h00;
  assign mem[1903] = 5'h01;
  assign mem[1904] = 5'h10;
  assign mem[1905] = 5'h00;
  assign mem[1906] = 5'h03;
  assign mem[1907] = 5'h12;
  assign mem[1908] = 5'h11;
  assign mem[1909] = 5'h10;
  assign mem[1910] = 5'h00;
  assign mem[1911] = 5'h01;
  assign mem[1912] = 5'h10;
  assign mem[1913] = 5'h00;
  assign mem[1914] = 5'h02;
  assign mem[1915] = 5'h11;
  assign mem[1916] = 5'h10;
  assign mem[1917] = 5'h00;
  assign mem[1918] = 5'h01;
  assign mem[1919] = 5'h10;
  assign mem[1920] = 5'h00;
  assign mem[1921] = 5'h06;
  assign mem[1922] = 5'h15;
  assign mem[1923] = 5'h14;
  assign mem[1924] = 5'h13;
  assign mem[1925] = 5'h12;
  assign mem[1926] = 5'h11;
  assign mem[1927] = 5'h10;
  assign mem[1928] = 5'h00;
  assign mem[1929] = 5'h01;
  assign mem[1930] = 5'h10;
  assign mem[1931] = 5'h00;
  assign mem[1932] = 5'h02;
  assign mem[1933] = 5'h11;
  assign mem[1934] = 5'h10;
  assign mem[1935] = 5'h00;
  assign mem[1936] = 5'h01;
  assign mem[1937] = 5'h10;
  assign mem[1938] = 5'h00;
  assign mem[1939] = 5'h03;
  assign mem[1940] = 5'h12;
  assign mem[1941] = 5'h11;
  assign mem[1942] = 5'h10;
  assign mem[1943] = 5'h00;
  assign mem[1944] = 5'h01;
  assign mem[1945] = 5'h10;
  assign mem[1946] = 5'h00;
  assign mem[1947] = 5'h02;
  assign mem[1948] = 5'h11;
  assign mem[1949] = 5'h10;
  assign mem[1950] = 5'h00;
  assign mem[1951] = 5'h01;
  assign mem[1952] = 5'h10;
  assign mem[1953] = 5'h00;
  assign mem[1954] = 5'h04;
  assign mem[1955] = 5'h13;
  assign mem[1956] = 5'h12;
  assign mem[1957] = 5'h11;
  assign mem[1958] = 5'h10;
  assign mem[1959] = 5'h00;
  assign mem[1960] = 5'h01;
  assign mem[1961] = 5'h10;
  assign mem[1962] = 5'h00;
  assign mem[1963] = 5'h02;
  assign mem[1964] = 5'h11;
  assign mem[1965] = 5'h10;
  assign mem[1966] = 5'h00;
  assign mem[1967] = 5'h01;
  assign mem[1968] = 5'h10;
  assign mem[1969] = 5'h00;
  assign mem[1970] = 5'h03;
  assign mem[1971] = 5'h12;
  assign mem[1972] = 5'h11;
  assign mem[1973] = 5'h10;
  assign mem[1974] = 5'h00;
  assign mem[1975] = 5'h01;
  assign mem[1976] = 5'h10;
  assign mem[1977] = 5'h00;
  assign mem[1978] = 5'h02;
  assign mem[1979] = 5'h11;
  assign mem[1980] = 5'h10;
  assign mem[1981] = 5'h00;
  assign mem[1982] = 5'h01;
  assign mem[1983] = 5'h10;
  assign mem[1984] = 5'h00;
  assign mem[1985] = 5'h05;
  assign mem[1986] = 5'h14;
  assign mem[1987] = 5'h13;
  assign mem[1988] = 5'h12;
  assign mem[1989] = 5'h11;
  assign mem[1990] = 5'h10;
  assign mem[1991] = 5'h00;
  assign mem[1992] = 5'h01;
  assign mem[1993] = 5'h10;
  assign mem[1994] = 5'h00;
  assign mem[1995] = 5'h02;
  assign mem[1996] = 5'h11;
  assign mem[1997] = 5'h10;
  assign mem[1998] = 5'h00;
  assign mem[1999] = 5'h01;
  assign mem[2000] = 5'h10;
  assign mem[2001] = 5'h00;
  assign mem[2002] = 5'h03;
  assign mem[2003] = 5'h12;
  assign mem[2004] = 5'h11;
  assign mem[2005] = 5'h10;
  assign mem[2006] = 5'h00;
  assign mem[2007] = 5'h01;
  assign mem[2008] = 5'h10;
  assign mem[2009] = 5'h00;
  assign mem[2010] = 5'h02;
  assign mem[2011] = 5'h11;
  assign mem[2012] = 5'h10;
  assign mem[2013] = 5'h00;
  assign mem[2014] = 5'h01;
  assign mem[2015] = 5'h10;
  assign mem[2016] = 5'h00;
  assign mem[2017] = 5'h04;
  assign mem[2018] = 5'h13;
  assign mem[2019] = 5'h12;
  assign mem[2020] = 5'h11;
  assign mem[2021] = 5'h10;
  assign mem[2022] = 5'h00;
  assign mem[2023] = 5'h01;
  assign mem[2024] = 5'h10;
  assign mem[2025] = 5'h00;
  assign mem[2026] = 5'h02;
  assign mem[2027] = 5'h11;
  assign mem[2028] = 5'h10;
  assign mem[2029] = 5'h00;
  assign mem[2030] = 5'h01;
  assign mem[2031] = 5'h10;
  assign mem[2032] = 5'h00;
  assign mem[2033] = 5'h03;
  assign mem[2034] = 5'h12;
  assign mem[2035] = 5'h11;
  assign mem[2036] = 5'h10;
  assign mem[2037] = 5'h00;
  assign mem[2038] = 5'h01;
  assign mem[2039] = 5'h10;
  assign mem[2040] = 5'h00;
  assign mem[2041] = 5'h02;
  assign mem[2042] = 5'h11;
  assign mem[2043] = 5'h10;
  assign mem[2044] = 5'h00;
  assign mem[2045] = 5'h01;
  assign mem[2046] = 5'h10;
  assign mem[2047] = 5'h00;
  assign mem[2048] = 5'h0a;
  assign mem[2049] = 5'h19;
  assign mem[2050] = 5'h18;
  assign mem[2051] = 5'h17;
  assign mem[2052] = 5'h16;
  assign mem[2053] = 5'h15;
  assign mem[2054] = 5'h14;
  assign mem[2055] = 5'h13;
  assign mem[2056] = 5'h12;
  assign mem[2057] = 5'h11;
  assign mem[2058] = 5'h10;
  assign mem[2059] = 5'h00;
  assign mem[2060] = 5'h01;
  assign mem[2061] = 5'h10;
  assign mem[2062] = 5'h00;
  assign mem[2063] = 5'h02;
  assign mem[2064] = 5'h11;
  assign mem[2065] = 5'h10;
  assign mem[2066] = 5'h00;
  assign mem[2067] = 5'h01;
  assign mem[2068] = 5'h10;
  assign mem[2069] = 5'h00;
  assign mem[2070] = 5'h03;
  assign mem[2071] = 5'h12;
  assign mem[2072] = 5'h11;
  assign mem[2073] = 5'h10;
  assign mem[2074] = 5'h00;
  assign mem[2075] = 5'h01;
  assign mem[2076] = 5'h10;
  assign mem[2077] = 5'h00;
  assign mem[2078] = 5'h02;
  assign mem[2079] = 5'h11;
  assign mem[2080] = 5'h10;
  assign mem[2081] = 5'h00;
  assign mem[2082] = 5'h01;
  assign mem[2083] = 5'h10;
  assign mem[2084] = 5'h00;
  assign mem[2085] = 5'h04;
  assign mem[2086] = 5'h13;
  assign mem[2087] = 5'h12;
  assign mem[2088] = 5'h11;
  assign mem[2089] = 5'h10;
  assign mem[2090] = 5'h00;
  assign mem[2091] = 5'h01;
  assign mem[2092] = 5'h10;
  assign mem[2093] = 5'h00;
  assign mem[2094] = 5'h02;
  assign mem[2095] = 5'h11;
  assign mem[2096] = 5'h10;
  assign mem[2097] = 5'h00;
  assign mem[2098] = 5'h01;
  assign mem[2099] = 5'h10;
  assign mem[2100] = 5'h00;
  assign mem[2101] = 5'h03;
  assign mem[2102] = 5'h12;
  assign mem[2103] = 5'h11;
  assign mem[2104] = 5'h10;
  assign mem[2105] = 5'h00;
  assign mem[2106] = 5'h01;
  assign mem[2107] = 5'h10;
  assign mem[2108] = 5'h00;
  assign mem[2109] = 5'h02;
  assign mem[2110] = 5'h11;
  assign mem[2111] = 5'h10;
  assign mem[2112] = 5'h00;
  assign mem[2113] = 5'h01;
  assign mem[2114] = 5'h10;
  assign mem[2115] = 5'h00;
  assign mem[2116] = 5'h05;
  assign mem[2117] = 5'h14;
  assign mem[2118] = 5'h13;
  assign mem[2119] = 5'h12;
  assign mem[2120] = 5'h11;
  assign mem[2121] = 5'h10;
  assign mem[2122] = 5'h00;
  assign mem[2123] = 5'h01;
  assign mem[2124] = 5'h10;
  assign mem[2125] = 5'h00;
  assign mem[2126] = 5'h02;
  assign mem[2127] = 5'h11;
  assign mem[2128] = 5'h10;
  assign mem[2129] = 5'h00;
  assign mem[2130] = 5'h01;
  assign mem[2131] = 5'h10;
  assign mem[2132] = 5'h00;
  assign mem[2133] = 5'h03;
  assign mem[2134] = 5'h12;
  assign mem[2135] = 5'h11;
  assign mem[2136] = 5'h10;
  assign mem[2137] = 5'h00;
  assign mem[2138] = 5'h01;
  assign mem[2139] = 5'h10;
  assign mem[2140] = 5'h00;
  assign mem[2141] = 5'h02;
  assign mem[2142] = 5'h11;
  assign mem[2143] = 5'h10;
  assign mem[2144] = 5'h00;
  assign mem[2145] = 5'h01;
  assign mem[2146] = 5'h10;
  assign mem[2147] = 5'h00;
  assign mem[2148] = 5'h04;
  assign mem[2149] = 5'h13;
  assign mem[2150] = 5'h12;
  assign mem[2151] = 5'h11;
  assign mem[2152] = 5'h10;
  assign mem[2153] = 5'h00;
  assign mem[2154] = 5'h01;
  assign mem[2155] = 5'h10;
  assign mem[2156] = 5'h00;
  assign mem[2157] = 5'h02;
  assign mem[2158] = 5'h11;
  assign mem[2159] = 5'h10;
  assign mem[2160] = 5'h00;
  assign mem[2161] = 5'h01;
  assign mem[2162] = 5'h10;
  assign mem[2163] = 5'h00;
  assign mem[2164] = 5'h03;
  assign mem[2165] = 5'h12;
  assign mem[2166] = 5'h11;
  assign mem[2167] = 5'h10;
  assign mem[2168] = 5'h00;
  assign mem[2169] = 5'h01;
  assign mem[2170] = 5'h10;
  assign mem[2171] = 5'h00;
  assign mem[2172] = 5'h02;
  assign mem[2173] = 5'h11;
  assign mem[2174] = 5'h10;
  assign mem[2175] = 5'h00;
  assign mem[2176] = 5'h01;
  assign mem[2177] = 5'h10;
  assign mem[2178] = 5'h00;
  assign mem[2179] = 5'h06;
  assign mem[2180] = 5'h15;
  assign mem[2181] = 5'h14;
  assign mem[2182] = 5'h13;
  assign mem[2183] = 5'h12;
  assign mem[2184] = 5'h11;
  assign mem[2185] = 5'h10;
  assign mem[2186] = 5'h00;
  assign mem[2187] = 5'h01;
  assign mem[2188] = 5'h10;
  assign mem[2189] = 5'h00;
  assign mem[2190] = 5'h02;
  assign mem[2191] = 5'h11;
  assign mem[2192] = 5'h10;
  assign mem[2193] = 5'h00;
  assign mem[2194] = 5'h01;
  assign mem[2195] = 5'h10;
  assign mem[2196] = 5'h00;
  assign mem[2197] = 5'h03;
  assign mem[2198] = 5'h12;
  assign mem[2199] = 5'h11;
  assign mem[2200] = 5'h10;
  assign mem[2201] = 5'h00;
  assign mem[2202] = 5'h01;
  assign mem[2203] = 5'h10;
  assign mem[2204] = 5'h00;
  assign mem[2205] = 5'h02;
  assign mem[2206] = 5'h11;
  assign mem[2207] = 5'h10;
  assign mem[2208] = 5'h00;
  assign mem[2209] = 5'h01;
  assign mem[2210] = 5'h10;
  assign mem[2211] = 5'h00;
  assign mem[2212] = 5'h04;
  assign mem[2213] = 5'h13;
  assign mem[2214] = 5'h12;
  assign mem[2215] = 5'h11;
  assign mem[2216] = 5'h10;
  assign mem[2217] = 5'h00;
  assign mem[2218] = 5'h01;
  assign mem[2219] = 5'h10;
  assign mem[2220] = 5'h00;
  assign mem[2221] = 5'h02;
  assign mem[2222] = 5'h11;
  assign mem[2223] = 5'h10;
  assign mem[2224] = 5'h00;
  assign mem[2225] = 5'h01;
  assign mem[2226] = 5'h10;
  assign mem[2227] = 5'h00;
  assign mem[2228] = 5'h03;
  assign mem[2229] = 5'h12;
  assign mem[2230] = 5'h11;
  assign mem[2231] = 5'h10;
  assign mem[2232] = 5'h00;
  assign mem[2233] = 5'h01;
  assign mem[2234] = 5'h10;
  assign mem[2235] = 5'h00;
  assign mem[2236] = 5'h02;
  assign mem[2237] = 5'h11;
  assign mem[2238] = 5'h10;
  assign mem[2239] = 5'h00;
  assign mem[2240] = 5'h01;
  assign mem[2241] = 5'h10;
  assign mem[2242] = 5'h00;
  assign mem[2243] = 5'h05;
  assign mem[2244] = 5'h14;
  assign mem[2245] = 5'h13;
  assign mem[2246] = 5'h12;
  assign mem[2247] = 5'h11;
  assign mem[2248] = 5'h10;
  assign mem[2249] = 5'h00;
  assign mem[2250] = 5'h01;
  assign mem[2251] = 5'h10;
  assign mem[2252] = 5'h00;
  assign mem[2253] = 5'h02;
  assign mem[2254] = 5'h11;
  assign mem[2255] = 5'h10;
  assign mem[2256] = 5'h00;
  assign mem[2257] = 5'h01;
  assign mem[2258] = 5'h10;
  assign mem[2259] = 5'h00;
  assign mem[2260] = 5'h03;
  assign mem[2261] = 5'h12;
  assign mem[2262] = 5'h11;
  assign mem[2263] = 5'h10;
  assign mem[2264] = 5'h00;
  assign mem[2265] = 5'h01;
  assign mem[2266] = 5'h10;
  assign mem[2267] = 5'h00;
  assign mem[2268] = 5'h02;
  assign mem[2269] = 5'h11;
  assign mem[2270] = 5'h10;
  assign mem[2271] = 5'h00;
  assign mem[2272] = 5'h01;
  assign mem[2273] = 5'h10;
  assign mem[2274] = 5'h00;
  assign mem[2275] = 5'h04;
  assign mem[2276] = 5'h13;
  assign mem[2277] = 5'h12;
  assign mem[2278] = 5'h11;
  assign mem[2279] = 5'h10;
  assign mem[2280] = 5'h00;
  assign mem[2281] = 5'h01;
  assign mem[2282] = 5'h10;
  assign mem[2283] = 5'h00;
  assign mem[2284] = 5'h02;
  assign mem[2285] = 5'h11;
  assign mem[2286] = 5'h10;
  assign mem[2287] = 5'h00;
  assign mem[2288] = 5'h01;
  assign mem[2289] = 5'h10;
  assign mem[2290] = 5'h00;
  assign mem[2291] = 5'h03;
  assign mem[2292] = 5'h12;
  assign mem[2293] = 5'h11;
  assign mem[2294] = 5'h10;
  assign mem[2295] = 5'h00;
  assign mem[2296] = 5'h01;
  assign mem[2297] = 5'h10;
  assign mem[2298] = 5'h00;
  assign mem[2299] = 5'h02;
  assign mem[2300] = 5'h11;
  assign mem[2301] = 5'h10;
  assign mem[2302] = 5'h00;
  assign mem[2303] = 5'h01;
  assign mem[2304] = 5'h10;
  assign mem[2305] = 5'h00;
  assign mem[2306] = 5'h07;
  assign mem[2307] = 5'h16;
  assign mem[2308] = 5'h15;
  assign mem[2309] = 5'h14;
  assign mem[2310] = 5'h13;
  assign mem[2311] = 5'h12;
  assign mem[2312] = 5'h11;
  assign mem[2313] = 5'h10;
  assign mem[2314] = 5'h00;
  assign mem[2315] = 5'h01;
  assign mem[2316] = 5'h10;
  assign mem[2317] = 5'h00;
  assign mem[2318] = 5'h02;
  assign mem[2319] = 5'h11;
  assign mem[2320] = 5'h10;
  assign mem[2321] = 5'h00;
  assign mem[2322] = 5'h01;
  assign mem[2323] = 5'h10;
  assign mem[2324] = 5'h00;
  assign mem[2325] = 5'h03;
  assign mem[2326] = 5'h12;
  assign mem[2327] = 5'h11;
  assign mem[2328] = 5'h10;
  assign mem[2329] = 5'h00;
  assign mem[2330] = 5'h01;
  assign mem[2331] = 5'h10;
  assign mem[2332] = 5'h00;
  assign mem[2333] = 5'h02;
  assign mem[2334] = 5'h11;
  assign mem[2335] = 5'h10;
  assign mem[2336] = 5'h00;
  assign mem[2337] = 5'h01;
  assign mem[2338] = 5'h10;
  assign mem[2339] = 5'h00;
  assign mem[2340] = 5'h04;
  assign mem[2341] = 5'h13;
  assign mem[2342] = 5'h12;
  assign mem[2343] = 5'h11;
  assign mem[2344] = 5'h10;
  assign mem[2345] = 5'h00;
  assign mem[2346] = 5'h01;
  assign mem[2347] = 5'h10;
  assign mem[2348] = 5'h00;
  assign mem[2349] = 5'h02;
  assign mem[2350] = 5'h11;
  assign mem[2351] = 5'h10;
  assign mem[2352] = 5'h00;
  assign mem[2353] = 5'h01;
  assign mem[2354] = 5'h10;
  assign mem[2355] = 5'h00;
  assign mem[2356] = 5'h03;
  assign mem[2357] = 5'h12;
  assign mem[2358] = 5'h11;
  assign mem[2359] = 5'h10;
  assign mem[2360] = 5'h00;
  assign mem[2361] = 5'h01;
  assign mem[2362] = 5'h10;
  assign mem[2363] = 5'h00;
  assign mem[2364] = 5'h02;
  assign mem[2365] = 5'h11;
  assign mem[2366] = 5'h10;
  assign mem[2367] = 5'h00;
  assign mem[2368] = 5'h01;
  assign mem[2369] = 5'h10;
  assign mem[2370] = 5'h00;
  assign mem[2371] = 5'h05;
  assign mem[2372] = 5'h14;
  assign mem[2373] = 5'h13;
  assign mem[2374] = 5'h12;
  assign mem[2375] = 5'h11;
  assign mem[2376] = 5'h10;
  assign mem[2377] = 5'h00;
  assign mem[2378] = 5'h01;
  assign mem[2379] = 5'h10;
  assign mem[2380] = 5'h00;
  assign mem[2381] = 5'h02;
  assign mem[2382] = 5'h11;
  assign mem[2383] = 5'h10;
  assign mem[2384] = 5'h00;
  assign mem[2385] = 5'h01;
  assign mem[2386] = 5'h10;
  assign mem[2387] = 5'h00;
  assign mem[2388] = 5'h03;
  assign mem[2389] = 5'h12;
  assign mem[2390] = 5'h11;
  assign mem[2391] = 5'h10;
  assign mem[2392] = 5'h00;
  assign mem[2393] = 5'h01;
  assign mem[2394] = 5'h10;
  assign mem[2395] = 5'h00;
  assign mem[2396] = 5'h02;
  assign mem[2397] = 5'h11;
  assign mem[2398] = 5'h10;
  assign mem[2399] = 5'h00;
  assign mem[2400] = 5'h01;
  assign mem[2401] = 5'h10;
  assign mem[2402] = 5'h00;
  assign mem[2403] = 5'h04;
  assign mem[2404] = 5'h13;
  assign mem[2405] = 5'h12;
  assign mem[2406] = 5'h11;
  assign mem[2407] = 5'h10;
  assign mem[2408] = 5'h00;
  assign mem[2409] = 5'h01;
  assign mem[2410] = 5'h10;
  assign mem[2411] = 5'h00;
  assign mem[2412] = 5'h02;
  assign mem[2413] = 5'h11;
  assign mem[2414] = 5'h10;
  assign mem[2415] = 5'h00;
  assign mem[2416] = 5'h01;
  assign mem[2417] = 5'h10;
  assign mem[2418] = 5'h00;
  assign mem[2419] = 5'h03;
  assign mem[2420] = 5'h12;
  assign mem[2421] = 5'h11;
  assign mem[2422] = 5'h10;
  assign mem[2423] = 5'h00;
  assign mem[2424] = 5'h01;
  assign mem[2425] = 5'h10;
  assign mem[2426] = 5'h00;
  assign mem[2427] = 5'h02;
  assign mem[2428] = 5'h11;
  assign mem[2429] = 5'h10;
  assign mem[2430] = 5'h00;
  assign mem[2431] = 5'h01;
  assign mem[2432] = 5'h10;
  assign mem[2433] = 5'h00;
  assign mem[2434] = 5'h06;
  assign mem[2435] = 5'h15;
  assign mem[2436] = 5'h14;
  assign mem[2437] = 5'h13;
  assign mem[2438] = 5'h12;
  assign mem[2439] = 5'h11;
  assign mem[2440] = 5'h10;
  assign mem[2441] = 5'h00;
  assign mem[2442] = 5'h01;
  assign mem[2443] = 5'h10;
  assign mem[2444] = 5'h00;
  assign mem[2445] = 5'h02;
  assign mem[2446] = 5'h11;
  assign mem[2447] = 5'h10;
  assign mem[2448] = 5'h00;
  assign mem[2449] = 5'h01;
  assign mem[2450] = 5'h10;
  assign mem[2451] = 5'h00;
  assign mem[2452] = 5'h03;
  assign mem[2453] = 5'h12;
  assign mem[2454] = 5'h11;
  assign mem[2455] = 5'h10;
  assign mem[2456] = 5'h00;
  assign mem[2457] = 5'h01;
  assign mem[2458] = 5'h10;
  assign mem[2459] = 5'h00;
  assign mem[2460] = 5'h02;
  assign mem[2461] = 5'h11;
  assign mem[2462] = 5'h10;
  assign mem[2463] = 5'h00;
  assign mem[2464] = 5'h01;
  assign mem[2465] = 5'h10;
  assign mem[2466] = 5'h00;
  assign mem[2467] = 5'h04;
  assign mem[2468] = 5'h13;
  assign mem[2469] = 5'h12;
  assign mem[2470] = 5'h11;
  assign mem[2471] = 5'h10;
  assign mem[2472] = 5'h00;
  assign mem[2473] = 5'h01;
  assign mem[2474] = 5'h10;
  assign mem[2475] = 5'h00;
  assign mem[2476] = 5'h02;
  assign mem[2477] = 5'h11;
  assign mem[2478] = 5'h10;
  assign mem[2479] = 5'h00;
  assign mem[2480] = 5'h01;
  assign mem[2481] = 5'h10;
  assign mem[2482] = 5'h00;
  assign mem[2483] = 5'h03;
  assign mem[2484] = 5'h12;
  assign mem[2485] = 5'h11;
  assign mem[2486] = 5'h10;
  assign mem[2487] = 5'h00;
  assign mem[2488] = 5'h01;
  assign mem[2489] = 5'h10;
  assign mem[2490] = 5'h00;
  assign mem[2491] = 5'h02;
  assign mem[2492] = 5'h11;
  assign mem[2493] = 5'h10;
  assign mem[2494] = 5'h00;
  assign mem[2495] = 5'h01;
  assign mem[2496] = 5'h10;
  assign mem[2497] = 5'h00;
  assign mem[2498] = 5'h05;
  assign mem[2499] = 5'h14;
  assign mem[2500] = 5'h13;
  assign mem[2501] = 5'h12;
  assign mem[2502] = 5'h11;
  assign mem[2503] = 5'h10;
  assign mem[2504] = 5'h00;
  assign mem[2505] = 5'h01;
  assign mem[2506] = 5'h10;
  assign mem[2507] = 5'h00;
  assign mem[2508] = 5'h02;
  assign mem[2509] = 5'h11;
  assign mem[2510] = 5'h10;
  assign mem[2511] = 5'h00;
  assign mem[2512] = 5'h01;
  assign mem[2513] = 5'h10;
  assign mem[2514] = 5'h00;
  assign mem[2515] = 5'h03;
  assign mem[2516] = 5'h12;
  assign mem[2517] = 5'h11;
  assign mem[2518] = 5'h10;
  assign mem[2519] = 5'h00;
  assign mem[2520] = 5'h01;
  assign mem[2521] = 5'h10;
  assign mem[2522] = 5'h00;
  assign mem[2523] = 5'h02;
  assign mem[2524] = 5'h11;
  assign mem[2525] = 5'h10;
  assign mem[2526] = 5'h00;
  assign mem[2527] = 5'h01;
  assign mem[2528] = 5'h10;
  assign mem[2529] = 5'h00;
  assign mem[2530] = 5'h04;
  assign mem[2531] = 5'h13;
  assign mem[2532] = 5'h12;
  assign mem[2533] = 5'h11;
  assign mem[2534] = 5'h10;
  assign mem[2535] = 5'h00;
  assign mem[2536] = 5'h01;
  assign mem[2537] = 5'h10;
  assign mem[2538] = 5'h00;
  assign mem[2539] = 5'h02;
  assign mem[2540] = 5'h11;
  assign mem[2541] = 5'h10;
  assign mem[2542] = 5'h00;
  assign mem[2543] = 5'h01;
  assign mem[2544] = 5'h10;
  assign mem[2545] = 5'h00;
  assign mem[2546] = 5'h03;
  assign mem[2547] = 5'h12;
  assign mem[2548] = 5'h11;
  assign mem[2549] = 5'h10;
  assign mem[2550] = 5'h00;
  assign mem[2551] = 5'h01;
  assign mem[2552] = 5'h10;
  assign mem[2553] = 5'h00;
  assign mem[2554] = 5'h02;
  assign mem[2555] = 5'h11;
  assign mem[2556] = 5'h10;
  assign mem[2557] = 5'h00;
  assign mem[2558] = 5'h01;
  assign mem[2559] = 5'h10;
  assign mem[2560] = 5'h00;
  assign mem[2561] = 5'h08;
  assign mem[2562] = 5'h17;
  assign mem[2563] = 5'h16;
  assign mem[2564] = 5'h15;
  assign mem[2565] = 5'h14;
  assign mem[2566] = 5'h13;
  assign mem[2567] = 5'h12;
  assign mem[2568] = 5'h11;
  assign mem[2569] = 5'h10;
  assign mem[2570] = 5'h00;
  assign mem[2571] = 5'h01;
  assign mem[2572] = 5'h10;
  assign mem[2573] = 5'h00;
  assign mem[2574] = 5'h02;
  assign mem[2575] = 5'h11;
  assign mem[2576] = 5'h10;
  assign mem[2577] = 5'h00;
  assign mem[2578] = 5'h01;
  assign mem[2579] = 5'h10;
  assign mem[2580] = 5'h00;
  assign mem[2581] = 5'h03;
  assign mem[2582] = 5'h12;
  assign mem[2583] = 5'h11;
  assign mem[2584] = 5'h10;
  assign mem[2585] = 5'h00;
  assign mem[2586] = 5'h01;
  assign mem[2587] = 5'h10;
  assign mem[2588] = 5'h00;
  assign mem[2589] = 5'h02;
  assign mem[2590] = 5'h11;
  assign mem[2591] = 5'h10;
  assign mem[2592] = 5'h00;
  assign mem[2593] = 5'h01;
  assign mem[2594] = 5'h10;
  assign mem[2595] = 5'h00;
  assign mem[2596] = 5'h04;
  assign mem[2597] = 5'h13;
  assign mem[2598] = 5'h12;
  assign mem[2599] = 5'h11;
  assign mem[2600] = 5'h10;
  assign mem[2601] = 5'h00;
  assign mem[2602] = 5'h01;
  assign mem[2603] = 5'h10;
  assign mem[2604] = 5'h00;
  assign mem[2605] = 5'h02;
  assign mem[2606] = 5'h11;
  assign mem[2607] = 5'h10;
  assign mem[2608] = 5'h00;
  assign mem[2609] = 5'h01;
  assign mem[2610] = 5'h10;
  assign mem[2611] = 5'h00;
  assign mem[2612] = 5'h03;
  assign mem[2613] = 5'h12;
  assign mem[2614] = 5'h11;
  assign mem[2615] = 5'h10;
  assign mem[2616] = 5'h00;
  assign mem[2617] = 5'h01;
  assign mem[2618] = 5'h10;
  assign mem[2619] = 5'h00;
  assign mem[2620] = 5'h02;
  assign mem[2621] = 5'h11;
  assign mem[2622] = 5'h10;
  assign mem[2623] = 5'h00;
  assign mem[2624] = 5'h01;
  assign mem[2625] = 5'h10;
  assign mem[2626] = 5'h00;
  assign mem[2627] = 5'h05;
  assign mem[2628] = 5'h14;
  assign mem[2629] = 5'h13;
  assign mem[2630] = 5'h12;
  assign mem[2631] = 5'h11;
  assign mem[2632] = 5'h10;
  assign mem[2633] = 5'h00;
  assign mem[2634] = 5'h01;
  assign mem[2635] = 5'h10;
  assign mem[2636] = 5'h00;
  assign mem[2637] = 5'h02;
  assign mem[2638] = 5'h11;
  assign mem[2639] = 5'h10;
  assign mem[2640] = 5'h00;
  assign mem[2641] = 5'h01;
  assign mem[2642] = 5'h10;
  assign mem[2643] = 5'h00;
  assign mem[2644] = 5'h03;
  assign mem[2645] = 5'h12;
  assign mem[2646] = 5'h11;
  assign mem[2647] = 5'h10;
  assign mem[2648] = 5'h00;
  assign mem[2649] = 5'h01;
  assign mem[2650] = 5'h10;
  assign mem[2651] = 5'h00;
  assign mem[2652] = 5'h02;
  assign mem[2653] = 5'h11;
  assign mem[2654] = 5'h10;
  assign mem[2655] = 5'h00;
  assign mem[2656] = 5'h01;
  assign mem[2657] = 5'h10;
  assign mem[2658] = 5'h00;
  assign mem[2659] = 5'h04;
  assign mem[2660] = 5'h13;
  assign mem[2661] = 5'h12;
  assign mem[2662] = 5'h11;
  assign mem[2663] = 5'h10;
  assign mem[2664] = 5'h00;
  assign mem[2665] = 5'h01;
  assign mem[2666] = 5'h10;
  assign mem[2667] = 5'h00;
  assign mem[2668] = 5'h02;
  assign mem[2669] = 5'h11;
  assign mem[2670] = 5'h10;
  assign mem[2671] = 5'h00;
  assign mem[2672] = 5'h01;
  assign mem[2673] = 5'h10;
  assign mem[2674] = 5'h00;
  assign mem[2675] = 5'h03;
  assign mem[2676] = 5'h12;
  assign mem[2677] = 5'h11;
  assign mem[2678] = 5'h10;
  assign mem[2679] = 5'h00;
  assign mem[2680] = 5'h01;
  assign mem[2681] = 5'h10;
  assign mem[2682] = 5'h00;
  assign mem[2683] = 5'h02;
  assign mem[2684] = 5'h11;
  assign mem[2685] = 5'h10;
  assign mem[2686] = 5'h00;
  assign mem[2687] = 5'h01;
  assign mem[2688] = 5'h10;
  assign mem[2689] = 5'h00;
  assign mem[2690] = 5'h06;
  assign mem[2691] = 5'h15;
  assign mem[2692] = 5'h14;
  assign mem[2693] = 5'h13;
  assign mem[2694] = 5'h12;
  assign mem[2695] = 5'h11;
  assign mem[2696] = 5'h10;
  assign mem[2697] = 5'h00;
  assign mem[2698] = 5'h01;
  assign mem[2699] = 5'h10;
  assign mem[2700] = 5'h00;
  assign mem[2701] = 5'h02;
  assign mem[2702] = 5'h11;
  assign mem[2703] = 5'h10;
  assign mem[2704] = 5'h00;
  assign mem[2705] = 5'h01;
  assign mem[2706] = 5'h10;
  assign mem[2707] = 5'h00;
  assign mem[2708] = 5'h03;
  assign mem[2709] = 5'h12;
  assign mem[2710] = 5'h11;
  assign mem[2711] = 5'h10;
  assign mem[2712] = 5'h00;
  assign mem[2713] = 5'h01;
  assign mem[2714] = 5'h10;
  assign mem[2715] = 5'h00;
  assign mem[2716] = 5'h02;
  assign mem[2717] = 5'h11;
  assign mem[2718] = 5'h10;
  assign mem[2719] = 5'h00;
  assign mem[2720] = 5'h01;
  assign mem[2721] = 5'h10;
  assign mem[2722] = 5'h00;
  assign mem[2723] = 5'h04;
  assign mem[2724] = 5'h13;
  assign mem[2725] = 5'h12;
  assign mem[2726] = 5'h11;
  assign mem[2727] = 5'h10;
  assign mem[2728] = 5'h00;
  assign mem[2729] = 5'h01;
  assign mem[2730] = 5'h10;
  assign mem[2731] = 5'h00;
  assign mem[2732] = 5'h02;
  assign mem[2733] = 5'h11;
  assign mem[2734] = 5'h10;
  assign mem[2735] = 5'h00;
  assign mem[2736] = 5'h01;
  assign mem[2737] = 5'h10;
  assign mem[2738] = 5'h00;
  assign mem[2739] = 5'h03;
  assign mem[2740] = 5'h12;
  assign mem[2741] = 5'h11;
  assign mem[2742] = 5'h10;
  assign mem[2743] = 5'h00;
  assign mem[2744] = 5'h01;
  assign mem[2745] = 5'h10;
  assign mem[2746] = 5'h00;
  assign mem[2747] = 5'h02;
  assign mem[2748] = 5'h11;
  assign mem[2749] = 5'h10;
  assign mem[2750] = 5'h00;
  assign mem[2751] = 5'h01;
  assign mem[2752] = 5'h10;
  assign mem[2753] = 5'h00;
  assign mem[2754] = 5'h05;
  assign mem[2755] = 5'h14;
  assign mem[2756] = 5'h13;
  assign mem[2757] = 5'h12;
  assign mem[2758] = 5'h11;
  assign mem[2759] = 5'h10;
  assign mem[2760] = 5'h00;
  assign mem[2761] = 5'h01;
  assign mem[2762] = 5'h10;
  assign mem[2763] = 5'h00;
  assign mem[2764] = 5'h02;
  assign mem[2765] = 5'h11;
  assign mem[2766] = 5'h10;
  assign mem[2767] = 5'h00;
  assign mem[2768] = 5'h01;
  assign mem[2769] = 5'h10;
  assign mem[2770] = 5'h00;
  assign mem[2771] = 5'h03;
  assign mem[2772] = 5'h12;
  assign mem[2773] = 5'h11;
  assign mem[2774] = 5'h10;
  assign mem[2775] = 5'h00;
  assign mem[2776] = 5'h01;
  assign mem[2777] = 5'h10;
  assign mem[2778] = 5'h00;
  assign mem[2779] = 5'h02;
  assign mem[2780] = 5'h11;
  assign mem[2781] = 5'h10;
  assign mem[2782] = 5'h00;
  assign mem[2783] = 5'h01;
  assign mem[2784] = 5'h10;
  assign mem[2785] = 5'h00;
  assign mem[2786] = 5'h04;
  assign mem[2787] = 5'h13;
  assign mem[2788] = 5'h12;
  assign mem[2789] = 5'h11;
  assign mem[2790] = 5'h10;
  assign mem[2791] = 5'h00;
  assign mem[2792] = 5'h01;
  assign mem[2793] = 5'h10;
  assign mem[2794] = 5'h00;
  assign mem[2795] = 5'h02;
  assign mem[2796] = 5'h11;
  assign mem[2797] = 5'h10;
  assign mem[2798] = 5'h00;
  assign mem[2799] = 5'h01;
  assign mem[2800] = 5'h10;
  assign mem[2801] = 5'h00;
  assign mem[2802] = 5'h03;
  assign mem[2803] = 5'h12;
  assign mem[2804] = 5'h11;
  assign mem[2805] = 5'h10;
  assign mem[2806] = 5'h00;
  assign mem[2807] = 5'h01;
  assign mem[2808] = 5'h10;
  assign mem[2809] = 5'h00;
  assign mem[2810] = 5'h02;
  assign mem[2811] = 5'h11;
  assign mem[2812] = 5'h10;
  assign mem[2813] = 5'h00;
  assign mem[2814] = 5'h01;
  assign mem[2815] = 5'h10;
  assign mem[2816] = 5'h00;
  assign mem[2817] = 5'h07;
  assign mem[2818] = 5'h16;
  assign mem[2819] = 5'h15;
  assign mem[2820] = 5'h14;
  assign mem[2821] = 5'h13;
  assign mem[2822] = 5'h12;
  assign mem[2823] = 5'h11;
  assign mem[2824] = 5'h10;
  assign mem[2825] = 5'h00;
  assign mem[2826] = 5'h01;
  assign mem[2827] = 5'h10;
  assign mem[2828] = 5'h00;
  assign mem[2829] = 5'h02;
  assign mem[2830] = 5'h11;
  assign mem[2831] = 5'h10;
  assign mem[2832] = 5'h00;
  assign mem[2833] = 5'h01;
  assign mem[2834] = 5'h10;
  assign mem[2835] = 5'h00;
  assign mem[2836] = 5'h03;
  assign mem[2837] = 5'h12;
  assign mem[2838] = 5'h11;
  assign mem[2839] = 5'h10;
  assign mem[2840] = 5'h00;
  assign mem[2841] = 5'h01;
  assign mem[2842] = 5'h10;
  assign mem[2843] = 5'h00;
  assign mem[2844] = 5'h02;
  assign mem[2845] = 5'h11;
  assign mem[2846] = 5'h10;
  assign mem[2847] = 5'h00;
  assign mem[2848] = 5'h01;
  assign mem[2849] = 5'h10;
  assign mem[2850] = 5'h00;
  assign mem[2851] = 5'h04;
  assign mem[2852] = 5'h13;
  assign mem[2853] = 5'h12;
  assign mem[2854] = 5'h11;
  assign mem[2855] = 5'h10;
  assign mem[2856] = 5'h00;
  assign mem[2857] = 5'h01;
  assign mem[2858] = 5'h10;
  assign mem[2859] = 5'h00;
  assign mem[2860] = 5'h02;
  assign mem[2861] = 5'h11;
  assign mem[2862] = 5'h10;
  assign mem[2863] = 5'h00;
  assign mem[2864] = 5'h01;
  assign mem[2865] = 5'h10;
  assign mem[2866] = 5'h00;
  assign mem[2867] = 5'h03;
  assign mem[2868] = 5'h12;
  assign mem[2869] = 5'h11;
  assign mem[2870] = 5'h10;
  assign mem[2871] = 5'h00;
  assign mem[2872] = 5'h01;
  assign mem[2873] = 5'h10;
  assign mem[2874] = 5'h00;
  assign mem[2875] = 5'h02;
  assign mem[2876] = 5'h11;
  assign mem[2877] = 5'h10;
  assign mem[2878] = 5'h00;
  assign mem[2879] = 5'h01;
  assign mem[2880] = 5'h10;
  assign mem[2881] = 5'h00;
  assign mem[2882] = 5'h05;
  assign mem[2883] = 5'h14;
  assign mem[2884] = 5'h13;
  assign mem[2885] = 5'h12;
  assign mem[2886] = 5'h11;
  assign mem[2887] = 5'h10;
  assign mem[2888] = 5'h00;
  assign mem[2889] = 5'h01;
  assign mem[2890] = 5'h10;
  assign mem[2891] = 5'h00;
  assign mem[2892] = 5'h02;
  assign mem[2893] = 5'h11;
  assign mem[2894] = 5'h10;
  assign mem[2895] = 5'h00;
  assign mem[2896] = 5'h01;
  assign mem[2897] = 5'h10;
  assign mem[2898] = 5'h00;
  assign mem[2899] = 5'h03;
  assign mem[2900] = 5'h12;
  assign mem[2901] = 5'h11;
  assign mem[2902] = 5'h10;
  assign mem[2903] = 5'h00;
  assign mem[2904] = 5'h01;
  assign mem[2905] = 5'h10;
  assign mem[2906] = 5'h00;
  assign mem[2907] = 5'h02;
  assign mem[2908] = 5'h11;
  assign mem[2909] = 5'h10;
  assign mem[2910] = 5'h00;
  assign mem[2911] = 5'h01;
  assign mem[2912] = 5'h10;
  assign mem[2913] = 5'h00;
  assign mem[2914] = 5'h04;
  assign mem[2915] = 5'h13;
  assign mem[2916] = 5'h12;
  assign mem[2917] = 5'h11;
  assign mem[2918] = 5'h10;
  assign mem[2919] = 5'h00;
  assign mem[2920] = 5'h01;
  assign mem[2921] = 5'h10;
  assign mem[2922] = 5'h00;
  assign mem[2923] = 5'h02;
  assign mem[2924] = 5'h11;
  assign mem[2925] = 5'h10;
  assign mem[2926] = 5'h00;
  assign mem[2927] = 5'h01;
  assign mem[2928] = 5'h10;
  assign mem[2929] = 5'h00;
  assign mem[2930] = 5'h03;
  assign mem[2931] = 5'h12;
  assign mem[2932] = 5'h11;
  assign mem[2933] = 5'h10;
  assign mem[2934] = 5'h00;
  assign mem[2935] = 5'h01;
  assign mem[2936] = 5'h10;
  assign mem[2937] = 5'h00;
  assign mem[2938] = 5'h02;
  assign mem[2939] = 5'h11;
  assign mem[2940] = 5'h10;
  assign mem[2941] = 5'h00;
  assign mem[2942] = 5'h01;
  assign mem[2943] = 5'h10;
  assign mem[2944] = 5'h00;
  assign mem[2945] = 5'h06;
  assign mem[2946] = 5'h15;
  assign mem[2947] = 5'h14;
  assign mem[2948] = 5'h13;
  assign mem[2949] = 5'h12;
  assign mem[2950] = 5'h11;
  assign mem[2951] = 5'h10;
  assign mem[2952] = 5'h00;
  assign mem[2953] = 5'h01;
  assign mem[2954] = 5'h10;
  assign mem[2955] = 5'h00;
  assign mem[2956] = 5'h02;
  assign mem[2957] = 5'h11;
  assign mem[2958] = 5'h10;
  assign mem[2959] = 5'h00;
  assign mem[2960] = 5'h01;
  assign mem[2961] = 5'h10;
  assign mem[2962] = 5'h00;
  assign mem[2963] = 5'h03;
  assign mem[2964] = 5'h12;
  assign mem[2965] = 5'h11;
  assign mem[2966] = 5'h10;
  assign mem[2967] = 5'h00;
  assign mem[2968] = 5'h01;
  assign mem[2969] = 5'h10;
  assign mem[2970] = 5'h00;
  assign mem[2971] = 5'h02;
  assign mem[2972] = 5'h11;
  assign mem[2973] = 5'h10;
  assign mem[2974] = 5'h00;
  assign mem[2975] = 5'h01;
  assign mem[2976] = 5'h10;
  assign mem[2977] = 5'h00;
  assign mem[2978] = 5'h04;
  assign mem[2979] = 5'h13;
  assign mem[2980] = 5'h12;
  assign mem[2981] = 5'h11;
  assign mem[2982] = 5'h10;
  assign mem[2983] = 5'h00;
  assign mem[2984] = 5'h01;
  assign mem[2985] = 5'h10;
  assign mem[2986] = 5'h00;
  assign mem[2987] = 5'h02;
  assign mem[2988] = 5'h11;
  assign mem[2989] = 5'h10;
  assign mem[2990] = 5'h00;
  assign mem[2991] = 5'h01;
  assign mem[2992] = 5'h10;
  assign mem[2993] = 5'h00;
  assign mem[2994] = 5'h03;
  assign mem[2995] = 5'h12;
  assign mem[2996] = 5'h11;
  assign mem[2997] = 5'h10;
  assign mem[2998] = 5'h00;
  assign mem[2999] = 5'h01;
  assign mem[3000] = 5'h10;
  assign mem[3001] = 5'h00;
  assign mem[3002] = 5'h02;
  assign mem[3003] = 5'h11;
  assign mem[3004] = 5'h10;
  assign mem[3005] = 5'h00;
  assign mem[3006] = 5'h01;
  assign mem[3007] = 5'h10;
  assign mem[3008] = 5'h00;
  assign mem[3009] = 5'h05;
  assign mem[3010] = 5'h14;
  assign mem[3011] = 5'h13;
  assign mem[3012] = 5'h12;
  assign mem[3013] = 5'h11;
  assign mem[3014] = 5'h10;
  assign mem[3015] = 5'h00;
  assign mem[3016] = 5'h01;
  assign mem[3017] = 5'h10;
  assign mem[3018] = 5'h00;
  assign mem[3019] = 5'h02;
  assign mem[3020] = 5'h11;
  assign mem[3021] = 5'h10;
  assign mem[3022] = 5'h00;
  assign mem[3023] = 5'h01;
  assign mem[3024] = 5'h10;
  assign mem[3025] = 5'h00;
  assign mem[3026] = 5'h03;
  assign mem[3027] = 5'h12;
  assign mem[3028] = 5'h11;
  assign mem[3029] = 5'h10;
  assign mem[3030] = 5'h00;
  assign mem[3031] = 5'h01;
  assign mem[3032] = 5'h10;
  assign mem[3033] = 5'h00;
  assign mem[3034] = 5'h02;
  assign mem[3035] = 5'h11;
  assign mem[3036] = 5'h10;
  assign mem[3037] = 5'h00;
  assign mem[3038] = 5'h01;
  assign mem[3039] = 5'h10;
  assign mem[3040] = 5'h00;
  assign mem[3041] = 5'h04;
  assign mem[3042] = 5'h13;
  assign mem[3043] = 5'h12;
  assign mem[3044] = 5'h11;
  assign mem[3045] = 5'h10;
  assign mem[3046] = 5'h00;
  assign mem[3047] = 5'h01;
  assign mem[3048] = 5'h10;
  assign mem[3049] = 5'h00;
  assign mem[3050] = 5'h02;
  assign mem[3051] = 5'h11;
  assign mem[3052] = 5'h10;
  assign mem[3053] = 5'h00;
  assign mem[3054] = 5'h01;
  assign mem[3055] = 5'h10;
  assign mem[3056] = 5'h00;
  assign mem[3057] = 5'h03;
  assign mem[3058] = 5'h12;
  assign mem[3059] = 5'h11;
  assign mem[3060] = 5'h10;
  assign mem[3061] = 5'h00;
  assign mem[3062] = 5'h01;
  assign mem[3063] = 5'h10;
  assign mem[3064] = 5'h00;
  assign mem[3065] = 5'h02;
  assign mem[3066] = 5'h11;
  assign mem[3067] = 5'h10;
  assign mem[3068] = 5'h00;
  assign mem[3069] = 5'h01;
  assign mem[3070] = 5'h10;
  assign mem[3071] = 5'h00;
  assign mem[3072] = 5'h09;
  assign mem[3073] = 5'h18;
  assign mem[3074] = 5'h17;
  assign mem[3075] = 5'h16;
  assign mem[3076] = 5'h15;
  assign mem[3077] = 5'h14;
  assign mem[3078] = 5'h13;
  assign mem[3079] = 5'h12;
  assign mem[3080] = 5'h11;
  assign mem[3081] = 5'h10;
  assign mem[3082] = 5'h00;
  assign mem[3083] = 5'h01;
  assign mem[3084] = 5'h10;
  assign mem[3085] = 5'h00;
  assign mem[3086] = 5'h02;
  assign mem[3087] = 5'h11;
  assign mem[3088] = 5'h10;
  assign mem[3089] = 5'h00;
  assign mem[3090] = 5'h01;
  assign mem[3091] = 5'h10;
  assign mem[3092] = 5'h00;
  assign mem[3093] = 5'h03;
  assign mem[3094] = 5'h12;
  assign mem[3095] = 5'h11;
  assign mem[3096] = 5'h10;
  assign mem[3097] = 5'h00;
  assign mem[3098] = 5'h01;
  assign mem[3099] = 5'h10;
  assign mem[3100] = 5'h00;
  assign mem[3101] = 5'h02;
  assign mem[3102] = 5'h11;
  assign mem[3103] = 5'h10;
  assign mem[3104] = 5'h00;
  assign mem[3105] = 5'h01;
  assign mem[3106] = 5'h10;
  assign mem[3107] = 5'h00;
  assign mem[3108] = 5'h04;
  assign mem[3109] = 5'h13;
  assign mem[3110] = 5'h12;
  assign mem[3111] = 5'h11;
  assign mem[3112] = 5'h10;
  assign mem[3113] = 5'h00;
  assign mem[3114] = 5'h01;
  assign mem[3115] = 5'h10;
  assign mem[3116] = 5'h00;
  assign mem[3117] = 5'h02;
  assign mem[3118] = 5'h11;
  assign mem[3119] = 5'h10;
  assign mem[3120] = 5'h00;
  assign mem[3121] = 5'h01;
  assign mem[3122] = 5'h10;
  assign mem[3123] = 5'h00;
  assign mem[3124] = 5'h03;
  assign mem[3125] = 5'h12;
  assign mem[3126] = 5'h11;
  assign mem[3127] = 5'h10;
  assign mem[3128] = 5'h00;
  assign mem[3129] = 5'h01;
  assign mem[3130] = 5'h10;
  assign mem[3131] = 5'h00;
  assign mem[3132] = 5'h02;
  assign mem[3133] = 5'h11;
  assign mem[3134] = 5'h10;
  assign mem[3135] = 5'h00;
  assign mem[3136] = 5'h01;
  assign mem[3137] = 5'h10;
  assign mem[3138] = 5'h00;
  assign mem[3139] = 5'h05;
  assign mem[3140] = 5'h14;
  assign mem[3141] = 5'h13;
  assign mem[3142] = 5'h12;
  assign mem[3143] = 5'h11;
  assign mem[3144] = 5'h10;
  assign mem[3145] = 5'h00;
  assign mem[3146] = 5'h01;
  assign mem[3147] = 5'h10;
  assign mem[3148] = 5'h00;
  assign mem[3149] = 5'h02;
  assign mem[3150] = 5'h11;
  assign mem[3151] = 5'h10;
  assign mem[3152] = 5'h00;
  assign mem[3153] = 5'h01;
  assign mem[3154] = 5'h10;
  assign mem[3155] = 5'h00;
  assign mem[3156] = 5'h03;
  assign mem[3157] = 5'h12;
  assign mem[3158] = 5'h11;
  assign mem[3159] = 5'h10;
  assign mem[3160] = 5'h00;
  assign mem[3161] = 5'h01;
  assign mem[3162] = 5'h10;
  assign mem[3163] = 5'h00;
  assign mem[3164] = 5'h02;
  assign mem[3165] = 5'h11;
  assign mem[3166] = 5'h10;
  assign mem[3167] = 5'h00;
  assign mem[3168] = 5'h01;
  assign mem[3169] = 5'h10;
  assign mem[3170] = 5'h00;
  assign mem[3171] = 5'h04;
  assign mem[3172] = 5'h13;
  assign mem[3173] = 5'h12;
  assign mem[3174] = 5'h11;
  assign mem[3175] = 5'h10;
  assign mem[3176] = 5'h00;
  assign mem[3177] = 5'h01;
  assign mem[3178] = 5'h10;
  assign mem[3179] = 5'h00;
  assign mem[3180] = 5'h02;
  assign mem[3181] = 5'h11;
  assign mem[3182] = 5'h10;
  assign mem[3183] = 5'h00;
  assign mem[3184] = 5'h01;
  assign mem[3185] = 5'h10;
  assign mem[3186] = 5'h00;
  assign mem[3187] = 5'h03;
  assign mem[3188] = 5'h12;
  assign mem[3189] = 5'h11;
  assign mem[3190] = 5'h10;
  assign mem[3191] = 5'h00;
  assign mem[3192] = 5'h01;
  assign mem[3193] = 5'h10;
  assign mem[3194] = 5'h00;
  assign mem[3195] = 5'h02;
  assign mem[3196] = 5'h11;
  assign mem[3197] = 5'h10;
  assign mem[3198] = 5'h00;
  assign mem[3199] = 5'h01;
  assign mem[3200] = 5'h10;
  assign mem[3201] = 5'h00;
  assign mem[3202] = 5'h06;
  assign mem[3203] = 5'h15;
  assign mem[3204] = 5'h14;
  assign mem[3205] = 5'h13;
  assign mem[3206] = 5'h12;
  assign mem[3207] = 5'h11;
  assign mem[3208] = 5'h10;
  assign mem[3209] = 5'h00;
  assign mem[3210] = 5'h01;
  assign mem[3211] = 5'h10;
  assign mem[3212] = 5'h00;
  assign mem[3213] = 5'h02;
  assign mem[3214] = 5'h11;
  assign mem[3215] = 5'h10;
  assign mem[3216] = 5'h00;
  assign mem[3217] = 5'h01;
  assign mem[3218] = 5'h10;
  assign mem[3219] = 5'h00;
  assign mem[3220] = 5'h03;
  assign mem[3221] = 5'h12;
  assign mem[3222] = 5'h11;
  assign mem[3223] = 5'h10;
  assign mem[3224] = 5'h00;
  assign mem[3225] = 5'h01;
  assign mem[3226] = 5'h10;
  assign mem[3227] = 5'h00;
  assign mem[3228] = 5'h02;
  assign mem[3229] = 5'h11;
  assign mem[3230] = 5'h10;
  assign mem[3231] = 5'h00;
  assign mem[3232] = 5'h01;
  assign mem[3233] = 5'h10;
  assign mem[3234] = 5'h00;
  assign mem[3235] = 5'h04;
  assign mem[3236] = 5'h13;
  assign mem[3237] = 5'h12;
  assign mem[3238] = 5'h11;
  assign mem[3239] = 5'h10;
  assign mem[3240] = 5'h00;
  assign mem[3241] = 5'h01;
  assign mem[3242] = 5'h10;
  assign mem[3243] = 5'h00;
  assign mem[3244] = 5'h02;
  assign mem[3245] = 5'h11;
  assign mem[3246] = 5'h10;
  assign mem[3247] = 5'h00;
  assign mem[3248] = 5'h01;
  assign mem[3249] = 5'h10;
  assign mem[3250] = 5'h00;
  assign mem[3251] = 5'h03;
  assign mem[3252] = 5'h12;
  assign mem[3253] = 5'h11;
  assign mem[3254] = 5'h10;
  assign mem[3255] = 5'h00;
  assign mem[3256] = 5'h01;
  assign mem[3257] = 5'h10;
  assign mem[3258] = 5'h00;
  assign mem[3259] = 5'h02;
  assign mem[3260] = 5'h11;
  assign mem[3261] = 5'h10;
  assign mem[3262] = 5'h00;
  assign mem[3263] = 5'h01;
  assign mem[3264] = 5'h10;
  assign mem[3265] = 5'h00;
  assign mem[3266] = 5'h05;
  assign mem[3267] = 5'h14;
  assign mem[3268] = 5'h13;
  assign mem[3269] = 5'h12;
  assign mem[3270] = 5'h11;
  assign mem[3271] = 5'h10;
  assign mem[3272] = 5'h00;
  assign mem[3273] = 5'h01;
  assign mem[3274] = 5'h10;
  assign mem[3275] = 5'h00;
  assign mem[3276] = 5'h02;
  assign mem[3277] = 5'h11;
  assign mem[3278] = 5'h10;
  assign mem[3279] = 5'h00;
  assign mem[3280] = 5'h01;
  assign mem[3281] = 5'h10;
  assign mem[3282] = 5'h00;
  assign mem[3283] = 5'h03;
  assign mem[3284] = 5'h12;
  assign mem[3285] = 5'h11;
  assign mem[3286] = 5'h10;
  assign mem[3287] = 5'h00;
  assign mem[3288] = 5'h01;
  assign mem[3289] = 5'h10;
  assign mem[3290] = 5'h00;
  assign mem[3291] = 5'h02;
  assign mem[3292] = 5'h11;
  assign mem[3293] = 5'h10;
  assign mem[3294] = 5'h00;
  assign mem[3295] = 5'h01;
  assign mem[3296] = 5'h10;
  assign mem[3297] = 5'h00;
  assign mem[3298] = 5'h04;
  assign mem[3299] = 5'h13;
  assign mem[3300] = 5'h12;
  assign mem[3301] = 5'h11;
  assign mem[3302] = 5'h10;
  assign mem[3303] = 5'h00;
  assign mem[3304] = 5'h01;
  assign mem[3305] = 5'h10;
  assign mem[3306] = 5'h00;
  assign mem[3307] = 5'h02;
  assign mem[3308] = 5'h11;
  assign mem[3309] = 5'h10;
  assign mem[3310] = 5'h00;
  assign mem[3311] = 5'h01;
  assign mem[3312] = 5'h10;
  assign mem[3313] = 5'h00;
  assign mem[3314] = 5'h03;
  assign mem[3315] = 5'h12;
  assign mem[3316] = 5'h11;
  assign mem[3317] = 5'h10;
  assign mem[3318] = 5'h00;
  assign mem[3319] = 5'h01;
  assign mem[3320] = 5'h10;
  assign mem[3321] = 5'h00;
  assign mem[3322] = 5'h02;
  assign mem[3323] = 5'h11;
  assign mem[3324] = 5'h10;
  assign mem[3325] = 5'h00;
  assign mem[3326] = 5'h01;
  assign mem[3327] = 5'h10;
  assign mem[3328] = 5'h00;
  assign mem[3329] = 5'h07;
  assign mem[3330] = 5'h16;
  assign mem[3331] = 5'h15;
  assign mem[3332] = 5'h14;
  assign mem[3333] = 5'h13;
  assign mem[3334] = 5'h12;
  assign mem[3335] = 5'h11;
  assign mem[3336] = 5'h10;
  assign mem[3337] = 5'h00;
  assign mem[3338] = 5'h01;
  assign mem[3339] = 5'h10;
  assign mem[3340] = 5'h00;
  assign mem[3341] = 5'h02;
  assign mem[3342] = 5'h11;
  assign mem[3343] = 5'h10;
  assign mem[3344] = 5'h00;
  assign mem[3345] = 5'h01;
  assign mem[3346] = 5'h10;
  assign mem[3347] = 5'h00;
  assign mem[3348] = 5'h03;
  assign mem[3349] = 5'h12;
  assign mem[3350] = 5'h11;
  assign mem[3351] = 5'h10;
  assign mem[3352] = 5'h00;
  assign mem[3353] = 5'h01;
  assign mem[3354] = 5'h10;
  assign mem[3355] = 5'h00;
  assign mem[3356] = 5'h02;
  assign mem[3357] = 5'h11;
  assign mem[3358] = 5'h10;
  assign mem[3359] = 5'h00;
  assign mem[3360] = 5'h01;
  assign mem[3361] = 5'h10;
  assign mem[3362] = 5'h00;
  assign mem[3363] = 5'h04;
  assign mem[3364] = 5'h13;
  assign mem[3365] = 5'h12;
  assign mem[3366] = 5'h11;
  assign mem[3367] = 5'h10;
  assign mem[3368] = 5'h00;
  assign mem[3369] = 5'h01;
  assign mem[3370] = 5'h10;
  assign mem[3371] = 5'h00;
  assign mem[3372] = 5'h02;
  assign mem[3373] = 5'h11;
  assign mem[3374] = 5'h10;
  assign mem[3375] = 5'h00;
  assign mem[3376] = 5'h01;
  assign mem[3377] = 5'h10;
  assign mem[3378] = 5'h00;
  assign mem[3379] = 5'h03;
  assign mem[3380] = 5'h12;
  assign mem[3381] = 5'h11;
  assign mem[3382] = 5'h10;
  assign mem[3383] = 5'h00;
  assign mem[3384] = 5'h01;
  assign mem[3385] = 5'h10;
  assign mem[3386] = 5'h00;
  assign mem[3387] = 5'h02;
  assign mem[3388] = 5'h11;
  assign mem[3389] = 5'h10;
  assign mem[3390] = 5'h00;
  assign mem[3391] = 5'h01;
  assign mem[3392] = 5'h10;
  assign mem[3393] = 5'h00;
  assign mem[3394] = 5'h05;
  assign mem[3395] = 5'h14;
  assign mem[3396] = 5'h13;
  assign mem[3397] = 5'h12;
  assign mem[3398] = 5'h11;
  assign mem[3399] = 5'h10;
  assign mem[3400] = 5'h00;
  assign mem[3401] = 5'h01;
  assign mem[3402] = 5'h10;
  assign mem[3403] = 5'h00;
  assign mem[3404] = 5'h02;
  assign mem[3405] = 5'h11;
  assign mem[3406] = 5'h10;
  assign mem[3407] = 5'h00;
  assign mem[3408] = 5'h01;
  assign mem[3409] = 5'h10;
  assign mem[3410] = 5'h00;
  assign mem[3411] = 5'h03;
  assign mem[3412] = 5'h12;
  assign mem[3413] = 5'h11;
  assign mem[3414] = 5'h10;
  assign mem[3415] = 5'h00;
  assign mem[3416] = 5'h01;
  assign mem[3417] = 5'h10;
  assign mem[3418] = 5'h00;
  assign mem[3419] = 5'h02;
  assign mem[3420] = 5'h11;
  assign mem[3421] = 5'h10;
  assign mem[3422] = 5'h00;
  assign mem[3423] = 5'h01;
  assign mem[3424] = 5'h10;
  assign mem[3425] = 5'h00;
  assign mem[3426] = 5'h04;
  assign mem[3427] = 5'h13;
  assign mem[3428] = 5'h12;
  assign mem[3429] = 5'h11;
  assign mem[3430] = 5'h10;
  assign mem[3431] = 5'h00;
  assign mem[3432] = 5'h01;
  assign mem[3433] = 5'h10;
  assign mem[3434] = 5'h00;
  assign mem[3435] = 5'h02;
  assign mem[3436] = 5'h11;
  assign mem[3437] = 5'h10;
  assign mem[3438] = 5'h00;
  assign mem[3439] = 5'h01;
  assign mem[3440] = 5'h10;
  assign mem[3441] = 5'h00;
  assign mem[3442] = 5'h03;
  assign mem[3443] = 5'h12;
  assign mem[3444] = 5'h11;
  assign mem[3445] = 5'h10;
  assign mem[3446] = 5'h00;
  assign mem[3447] = 5'h01;
  assign mem[3448] = 5'h10;
  assign mem[3449] = 5'h00;
  assign mem[3450] = 5'h02;
  assign mem[3451] = 5'h11;
  assign mem[3452] = 5'h10;
  assign mem[3453] = 5'h00;
  assign mem[3454] = 5'h01;
  assign mem[3455] = 5'h10;
  assign mem[3456] = 5'h00;
  assign mem[3457] = 5'h06;
  assign mem[3458] = 5'h15;
  assign mem[3459] = 5'h14;
  assign mem[3460] = 5'h13;
  assign mem[3461] = 5'h12;
  assign mem[3462] = 5'h11;
  assign mem[3463] = 5'h10;
  assign mem[3464] = 5'h00;
  assign mem[3465] = 5'h01;
  assign mem[3466] = 5'h10;
  assign mem[3467] = 5'h00;
  assign mem[3468] = 5'h02;
  assign mem[3469] = 5'h11;
  assign mem[3470] = 5'h10;
  assign mem[3471] = 5'h00;
  assign mem[3472] = 5'h01;
  assign mem[3473] = 5'h10;
  assign mem[3474] = 5'h00;
  assign mem[3475] = 5'h03;
  assign mem[3476] = 5'h12;
  assign mem[3477] = 5'h11;
  assign mem[3478] = 5'h10;
  assign mem[3479] = 5'h00;
  assign mem[3480] = 5'h01;
  assign mem[3481] = 5'h10;
  assign mem[3482] = 5'h00;
  assign mem[3483] = 5'h02;
  assign mem[3484] = 5'h11;
  assign mem[3485] = 5'h10;
  assign mem[3486] = 5'h00;
  assign mem[3487] = 5'h01;
  assign mem[3488] = 5'h10;
  assign mem[3489] = 5'h00;
  assign mem[3490] = 5'h04;
  assign mem[3491] = 5'h13;
  assign mem[3492] = 5'h12;
  assign mem[3493] = 5'h11;
  assign mem[3494] = 5'h10;
  assign mem[3495] = 5'h00;
  assign mem[3496] = 5'h01;
  assign mem[3497] = 5'h10;
  assign mem[3498] = 5'h00;
  assign mem[3499] = 5'h02;
  assign mem[3500] = 5'h11;
  assign mem[3501] = 5'h10;
  assign mem[3502] = 5'h00;
  assign mem[3503] = 5'h01;
  assign mem[3504] = 5'h10;
  assign mem[3505] = 5'h00;
  assign mem[3506] = 5'h03;
  assign mem[3507] = 5'h12;
  assign mem[3508] = 5'h11;
  assign mem[3509] = 5'h10;
  assign mem[3510] = 5'h00;
  assign mem[3511] = 5'h01;
  assign mem[3512] = 5'h10;
  assign mem[3513] = 5'h00;
  assign mem[3514] = 5'h02;
  assign mem[3515] = 5'h11;
  assign mem[3516] = 5'h10;
  assign mem[3517] = 5'h00;
  assign mem[3518] = 5'h01;
  assign mem[3519] = 5'h10;
  assign mem[3520] = 5'h00;
  assign mem[3521] = 5'h05;
  assign mem[3522] = 5'h14;
  assign mem[3523] = 5'h13;
  assign mem[3524] = 5'h12;
  assign mem[3525] = 5'h11;
  assign mem[3526] = 5'h10;
  assign mem[3527] = 5'h00;
  assign mem[3528] = 5'h01;
  assign mem[3529] = 5'h10;
  assign mem[3530] = 5'h00;
  assign mem[3531] = 5'h02;
  assign mem[3532] = 5'h11;
  assign mem[3533] = 5'h10;
  assign mem[3534] = 5'h00;
  assign mem[3535] = 5'h01;
  assign mem[3536] = 5'h10;
  assign mem[3537] = 5'h00;
  assign mem[3538] = 5'h03;
  assign mem[3539] = 5'h12;
  assign mem[3540] = 5'h11;
  assign mem[3541] = 5'h10;
  assign mem[3542] = 5'h00;
  assign mem[3543] = 5'h01;
  assign mem[3544] = 5'h10;
  assign mem[3545] = 5'h00;
  assign mem[3546] = 5'h02;
  assign mem[3547] = 5'h11;
  assign mem[3548] = 5'h10;
  assign mem[3549] = 5'h00;
  assign mem[3550] = 5'h01;
  assign mem[3551] = 5'h10;
  assign mem[3552] = 5'h00;
  assign mem[3553] = 5'h04;
  assign mem[3554] = 5'h13;
  assign mem[3555] = 5'h12;
  assign mem[3556] = 5'h11;
  assign mem[3557] = 5'h10;
  assign mem[3558] = 5'h00;
  assign mem[3559] = 5'h01;
  assign mem[3560] = 5'h10;
  assign mem[3561] = 5'h00;
  assign mem[3562] = 5'h02;
  assign mem[3563] = 5'h11;
  assign mem[3564] = 5'h10;
  assign mem[3565] = 5'h00;
  assign mem[3566] = 5'h01;
  assign mem[3567] = 5'h10;
  assign mem[3568] = 5'h00;
  assign mem[3569] = 5'h03;
  assign mem[3570] = 5'h12;
  assign mem[3571] = 5'h11;
  assign mem[3572] = 5'h10;
  assign mem[3573] = 5'h00;
  assign mem[3574] = 5'h01;
  assign mem[3575] = 5'h10;
  assign mem[3576] = 5'h00;
  assign mem[3577] = 5'h02;
  assign mem[3578] = 5'h11;
  assign mem[3579] = 5'h10;
  assign mem[3580] = 5'h00;
  assign mem[3581] = 5'h01;
  assign mem[3582] = 5'h10;
  assign mem[3583] = 5'h00;
  assign mem[3584] = 5'h08;
  assign mem[3585] = 5'h17;
  assign mem[3586] = 5'h16;
  assign mem[3587] = 5'h15;
  assign mem[3588] = 5'h14;
  assign mem[3589] = 5'h13;
  assign mem[3590] = 5'h12;
  assign mem[3591] = 5'h11;
  assign mem[3592] = 5'h10;
  assign mem[3593] = 5'h00;
  assign mem[3594] = 5'h01;
  assign mem[3595] = 5'h10;
  assign mem[3596] = 5'h00;
  assign mem[3597] = 5'h02;
  assign mem[3598] = 5'h11;
  assign mem[3599] = 5'h10;
  assign mem[3600] = 5'h00;
  assign mem[3601] = 5'h01;
  assign mem[3602] = 5'h10;
  assign mem[3603] = 5'h00;
  assign mem[3604] = 5'h03;
  assign mem[3605] = 5'h12;
  assign mem[3606] = 5'h11;
  assign mem[3607] = 5'h10;
  assign mem[3608] = 5'h00;
  assign mem[3609] = 5'h01;
  assign mem[3610] = 5'h10;
  assign mem[3611] = 5'h00;
  assign mem[3612] = 5'h02;
  assign mem[3613] = 5'h11;
  assign mem[3614] = 5'h10;
  assign mem[3615] = 5'h00;
  assign mem[3616] = 5'h01;
  assign mem[3617] = 5'h10;
  assign mem[3618] = 5'h00;
  assign mem[3619] = 5'h04;
  assign mem[3620] = 5'h13;
  assign mem[3621] = 5'h12;
  assign mem[3622] = 5'h11;
  assign mem[3623] = 5'h10;
  assign mem[3624] = 5'h00;
  assign mem[3625] = 5'h01;
  assign mem[3626] = 5'h10;
  assign mem[3627] = 5'h00;
  assign mem[3628] = 5'h02;
  assign mem[3629] = 5'h11;
  assign mem[3630] = 5'h10;
  assign mem[3631] = 5'h00;
  assign mem[3632] = 5'h01;
  assign mem[3633] = 5'h10;
  assign mem[3634] = 5'h00;
  assign mem[3635] = 5'h03;
  assign mem[3636] = 5'h12;
  assign mem[3637] = 5'h11;
  assign mem[3638] = 5'h10;
  assign mem[3639] = 5'h00;
  assign mem[3640] = 5'h01;
  assign mem[3641] = 5'h10;
  assign mem[3642] = 5'h00;
  assign mem[3643] = 5'h02;
  assign mem[3644] = 5'h11;
  assign mem[3645] = 5'h10;
  assign mem[3646] = 5'h00;
  assign mem[3647] = 5'h01;
  assign mem[3648] = 5'h10;
  assign mem[3649] = 5'h00;
  assign mem[3650] = 5'h05;
  assign mem[3651] = 5'h14;
  assign mem[3652] = 5'h13;
  assign mem[3653] = 5'h12;
  assign mem[3654] = 5'h11;
  assign mem[3655] = 5'h10;
  assign mem[3656] = 5'h00;
  assign mem[3657] = 5'h01;
  assign mem[3658] = 5'h10;
  assign mem[3659] = 5'h00;
  assign mem[3660] = 5'h02;
  assign mem[3661] = 5'h11;
  assign mem[3662] = 5'h10;
  assign mem[3663] = 5'h00;
  assign mem[3664] = 5'h01;
  assign mem[3665] = 5'h10;
  assign mem[3666] = 5'h00;
  assign mem[3667] = 5'h03;
  assign mem[3668] = 5'h12;
  assign mem[3669] = 5'h11;
  assign mem[3670] = 5'h10;
  assign mem[3671] = 5'h00;
  assign mem[3672] = 5'h01;
  assign mem[3673] = 5'h10;
  assign mem[3674] = 5'h00;
  assign mem[3675] = 5'h02;
  assign mem[3676] = 5'h11;
  assign mem[3677] = 5'h10;
  assign mem[3678] = 5'h00;
  assign mem[3679] = 5'h01;
  assign mem[3680] = 5'h10;
  assign mem[3681] = 5'h00;
  assign mem[3682] = 5'h04;
  assign mem[3683] = 5'h13;
  assign mem[3684] = 5'h12;
  assign mem[3685] = 5'h11;
  assign mem[3686] = 5'h10;
  assign mem[3687] = 5'h00;
  assign mem[3688] = 5'h01;
  assign mem[3689] = 5'h10;
  assign mem[3690] = 5'h00;
  assign mem[3691] = 5'h02;
  assign mem[3692] = 5'h11;
  assign mem[3693] = 5'h10;
  assign mem[3694] = 5'h00;
  assign mem[3695] = 5'h01;
  assign mem[3696] = 5'h10;
  assign mem[3697] = 5'h00;
  assign mem[3698] = 5'h03;
  assign mem[3699] = 5'h12;
  assign mem[3700] = 5'h11;
  assign mem[3701] = 5'h10;
  assign mem[3702] = 5'h00;
  assign mem[3703] = 5'h01;
  assign mem[3704] = 5'h10;
  assign mem[3705] = 5'h00;
  assign mem[3706] = 5'h02;
  assign mem[3707] = 5'h11;
  assign mem[3708] = 5'h10;
  assign mem[3709] = 5'h00;
  assign mem[3710] = 5'h01;
  assign mem[3711] = 5'h10;
  assign mem[3712] = 5'h00;
  assign mem[3713] = 5'h06;
  assign mem[3714] = 5'h15;
  assign mem[3715] = 5'h14;
  assign mem[3716] = 5'h13;
  assign mem[3717] = 5'h12;
  assign mem[3718] = 5'h11;
  assign mem[3719] = 5'h10;
  assign mem[3720] = 5'h00;
  assign mem[3721] = 5'h01;
  assign mem[3722] = 5'h10;
  assign mem[3723] = 5'h00;
  assign mem[3724] = 5'h02;
  assign mem[3725] = 5'h11;
  assign mem[3726] = 5'h10;
  assign mem[3727] = 5'h00;
  assign mem[3728] = 5'h01;
  assign mem[3729] = 5'h10;
  assign mem[3730] = 5'h00;
  assign mem[3731] = 5'h03;
  assign mem[3732] = 5'h12;
  assign mem[3733] = 5'h11;
  assign mem[3734] = 5'h10;
  assign mem[3735] = 5'h00;
  assign mem[3736] = 5'h01;
  assign mem[3737] = 5'h10;
  assign mem[3738] = 5'h00;
  assign mem[3739] = 5'h02;
  assign mem[3740] = 5'h11;
  assign mem[3741] = 5'h10;
  assign mem[3742] = 5'h00;
  assign mem[3743] = 5'h01;
  assign mem[3744] = 5'h10;
  assign mem[3745] = 5'h00;
  assign mem[3746] = 5'h04;
  assign mem[3747] = 5'h13;
  assign mem[3748] = 5'h12;
  assign mem[3749] = 5'h11;
  assign mem[3750] = 5'h10;
  assign mem[3751] = 5'h00;
  assign mem[3752] = 5'h01;
  assign mem[3753] = 5'h10;
  assign mem[3754] = 5'h00;
  assign mem[3755] = 5'h02;
  assign mem[3756] = 5'h11;
  assign mem[3757] = 5'h10;
  assign mem[3758] = 5'h00;
  assign mem[3759] = 5'h01;
  assign mem[3760] = 5'h10;
  assign mem[3761] = 5'h00;
  assign mem[3762] = 5'h03;
  assign mem[3763] = 5'h12;
  assign mem[3764] = 5'h11;
  assign mem[3765] = 5'h10;
  assign mem[3766] = 5'h00;
  assign mem[3767] = 5'h01;
  assign mem[3768] = 5'h10;
  assign mem[3769] = 5'h00;
  assign mem[3770] = 5'h02;
  assign mem[3771] = 5'h11;
  assign mem[3772] = 5'h10;
  assign mem[3773] = 5'h00;
  assign mem[3774] = 5'h01;
  assign mem[3775] = 5'h10;
  assign mem[3776] = 5'h00;
  assign mem[3777] = 5'h05;
  assign mem[3778] = 5'h14;
  assign mem[3779] = 5'h13;
  assign mem[3780] = 5'h12;
  assign mem[3781] = 5'h11;
  assign mem[3782] = 5'h10;
  assign mem[3783] = 5'h00;
  assign mem[3784] = 5'h01;
  assign mem[3785] = 5'h10;
  assign mem[3786] = 5'h00;
  assign mem[3787] = 5'h02;
  assign mem[3788] = 5'h11;
  assign mem[3789] = 5'h10;
  assign mem[3790] = 5'h00;
  assign mem[3791] = 5'h01;
  assign mem[3792] = 5'h10;
  assign mem[3793] = 5'h00;
  assign mem[3794] = 5'h03;
  assign mem[3795] = 5'h12;
  assign mem[3796] = 5'h11;
  assign mem[3797] = 5'h10;
  assign mem[3798] = 5'h00;
  assign mem[3799] = 5'h01;
  assign mem[3800] = 5'h10;
  assign mem[3801] = 5'h00;
  assign mem[3802] = 5'h02;
  assign mem[3803] = 5'h11;
  assign mem[3804] = 5'h10;
  assign mem[3805] = 5'h00;
  assign mem[3806] = 5'h01;
  assign mem[3807] = 5'h10;
  assign mem[3808] = 5'h00;
  assign mem[3809] = 5'h04;
  assign mem[3810] = 5'h13;
  assign mem[3811] = 5'h12;
  assign mem[3812] = 5'h11;
  assign mem[3813] = 5'h10;
  assign mem[3814] = 5'h00;
  assign mem[3815] = 5'h01;
  assign mem[3816] = 5'h10;
  assign mem[3817] = 5'h00;
  assign mem[3818] = 5'h02;
  assign mem[3819] = 5'h11;
  assign mem[3820] = 5'h10;
  assign mem[3821] = 5'h00;
  assign mem[3822] = 5'h01;
  assign mem[3823] = 5'h10;
  assign mem[3824] = 5'h00;
  assign mem[3825] = 5'h03;
  assign mem[3826] = 5'h12;
  assign mem[3827] = 5'h11;
  assign mem[3828] = 5'h10;
  assign mem[3829] = 5'h00;
  assign mem[3830] = 5'h01;
  assign mem[3831] = 5'h10;
  assign mem[3832] = 5'h00;
  assign mem[3833] = 5'h02;
  assign mem[3834] = 5'h11;
  assign mem[3835] = 5'h10;
  assign mem[3836] = 5'h00;
  assign mem[3837] = 5'h01;
  assign mem[3838] = 5'h10;
  assign mem[3839] = 5'h00;
  assign mem[3840] = 5'h07;
  assign mem[3841] = 5'h16;
  assign mem[3842] = 5'h15;
  assign mem[3843] = 5'h14;
  assign mem[3844] = 5'h13;
  assign mem[3845] = 5'h12;
  assign mem[3846] = 5'h11;
  assign mem[3847] = 5'h10;
  assign mem[3848] = 5'h00;
  assign mem[3849] = 5'h01;
  assign mem[3850] = 5'h10;
  assign mem[3851] = 5'h00;
  assign mem[3852] = 5'h02;
  assign mem[3853] = 5'h11;
  assign mem[3854] = 5'h10;
  assign mem[3855] = 5'h00;
  assign mem[3856] = 5'h01;
  assign mem[3857] = 5'h10;
  assign mem[3858] = 5'h00;
  assign mem[3859] = 5'h03;
  assign mem[3860] = 5'h12;
  assign mem[3861] = 5'h11;
  assign mem[3862] = 5'h10;
  assign mem[3863] = 5'h00;
  assign mem[3864] = 5'h01;
  assign mem[3865] = 5'h10;
  assign mem[3866] = 5'h00;
  assign mem[3867] = 5'h02;
  assign mem[3868] = 5'h11;
  assign mem[3869] = 5'h10;
  assign mem[3870] = 5'h00;
  assign mem[3871] = 5'h01;
  assign mem[3872] = 5'h10;
  assign mem[3873] = 5'h00;
  assign mem[3874] = 5'h04;
  assign mem[3875] = 5'h13;
  assign mem[3876] = 5'h12;
  assign mem[3877] = 5'h11;
  assign mem[3878] = 5'h10;
  assign mem[3879] = 5'h00;
  assign mem[3880] = 5'h01;
  assign mem[3881] = 5'h10;
  assign mem[3882] = 5'h00;
  assign mem[3883] = 5'h02;
  assign mem[3884] = 5'h11;
  assign mem[3885] = 5'h10;
  assign mem[3886] = 5'h00;
  assign mem[3887] = 5'h01;
  assign mem[3888] = 5'h10;
  assign mem[3889] = 5'h00;
  assign mem[3890] = 5'h03;
  assign mem[3891] = 5'h12;
  assign mem[3892] = 5'h11;
  assign mem[3893] = 5'h10;
  assign mem[3894] = 5'h00;
  assign mem[3895] = 5'h01;
  assign mem[3896] = 5'h10;
  assign mem[3897] = 5'h00;
  assign mem[3898] = 5'h02;
  assign mem[3899] = 5'h11;
  assign mem[3900] = 5'h10;
  assign mem[3901] = 5'h00;
  assign mem[3902] = 5'h01;
  assign mem[3903] = 5'h10;
  assign mem[3904] = 5'h00;
  assign mem[3905] = 5'h05;
  assign mem[3906] = 5'h14;
  assign mem[3907] = 5'h13;
  assign mem[3908] = 5'h12;
  assign mem[3909] = 5'h11;
  assign mem[3910] = 5'h10;
  assign mem[3911] = 5'h00;
  assign mem[3912] = 5'h01;
  assign mem[3913] = 5'h10;
  assign mem[3914] = 5'h00;
  assign mem[3915] = 5'h02;
  assign mem[3916] = 5'h11;
  assign mem[3917] = 5'h10;
  assign mem[3918] = 5'h00;
  assign mem[3919] = 5'h01;
  assign mem[3920] = 5'h10;
  assign mem[3921] = 5'h00;
  assign mem[3922] = 5'h03;
  assign mem[3923] = 5'h12;
  assign mem[3924] = 5'h11;
  assign mem[3925] = 5'h10;
  assign mem[3926] = 5'h00;
  assign mem[3927] = 5'h01;
  assign mem[3928] = 5'h10;
  assign mem[3929] = 5'h00;
  assign mem[3930] = 5'h02;
  assign mem[3931] = 5'h11;
  assign mem[3932] = 5'h10;
  assign mem[3933] = 5'h00;
  assign mem[3934] = 5'h01;
  assign mem[3935] = 5'h10;
  assign mem[3936] = 5'h00;
  assign mem[3937] = 5'h04;
  assign mem[3938] = 5'h13;
  assign mem[3939] = 5'h12;
  assign mem[3940] = 5'h11;
  assign mem[3941] = 5'h10;
  assign mem[3942] = 5'h00;
  assign mem[3943] = 5'h01;
  assign mem[3944] = 5'h10;
  assign mem[3945] = 5'h00;
  assign mem[3946] = 5'h02;
  assign mem[3947] = 5'h11;
  assign mem[3948] = 5'h10;
  assign mem[3949] = 5'h00;
  assign mem[3950] = 5'h01;
  assign mem[3951] = 5'h10;
  assign mem[3952] = 5'h00;
  assign mem[3953] = 5'h03;
  assign mem[3954] = 5'h12;
  assign mem[3955] = 5'h11;
  assign mem[3956] = 5'h10;
  assign mem[3957] = 5'h00;
  assign mem[3958] = 5'h01;
  assign mem[3959] = 5'h10;
  assign mem[3960] = 5'h00;
  assign mem[3961] = 5'h02;
  assign mem[3962] = 5'h11;
  assign mem[3963] = 5'h10;
  assign mem[3964] = 5'h00;
  assign mem[3965] = 5'h01;
  assign mem[3966] = 5'h10;
  assign mem[3967] = 5'h00;
  assign mem[3968] = 5'h06;
  assign mem[3969] = 5'h15;
  assign mem[3970] = 5'h14;
  assign mem[3971] = 5'h13;
  assign mem[3972] = 5'h12;
  assign mem[3973] = 5'h11;
  assign mem[3974] = 5'h10;
  assign mem[3975] = 5'h00;
  assign mem[3976] = 5'h01;
  assign mem[3977] = 5'h10;
  assign mem[3978] = 5'h00;
  assign mem[3979] = 5'h02;
  assign mem[3980] = 5'h11;
  assign mem[3981] = 5'h10;
  assign mem[3982] = 5'h00;
  assign mem[3983] = 5'h01;
  assign mem[3984] = 5'h10;
  assign mem[3985] = 5'h00;
  assign mem[3986] = 5'h03;
  assign mem[3987] = 5'h12;
  assign mem[3988] = 5'h11;
  assign mem[3989] = 5'h10;
  assign mem[3990] = 5'h00;
  assign mem[3991] = 5'h01;
  assign mem[3992] = 5'h10;
  assign mem[3993] = 5'h00;
  assign mem[3994] = 5'h02;
  assign mem[3995] = 5'h11;
  assign mem[3996] = 5'h10;
  assign mem[3997] = 5'h00;
  assign mem[3998] = 5'h01;
  assign mem[3999] = 5'h10;
  assign mem[4000] = 5'h00;
  assign mem[4001] = 5'h04;
  assign mem[4002] = 5'h13;
  assign mem[4003] = 5'h12;
  assign mem[4004] = 5'h11;
  assign mem[4005] = 5'h10;
  assign mem[4006] = 5'h00;
  assign mem[4007] = 5'h01;
  assign mem[4008] = 5'h10;
  assign mem[4009] = 5'h00;
  assign mem[4010] = 5'h02;
  assign mem[4011] = 5'h11;
  assign mem[4012] = 5'h10;
  assign mem[4013] = 5'h00;
  assign mem[4014] = 5'h01;
  assign mem[4015] = 5'h10;
  assign mem[4016] = 5'h00;
  assign mem[4017] = 5'h03;
  assign mem[4018] = 5'h12;
  assign mem[4019] = 5'h11;
  assign mem[4020] = 5'h10;
  assign mem[4021] = 5'h00;
  assign mem[4022] = 5'h01;
  assign mem[4023] = 5'h10;
  assign mem[4024] = 5'h00;
  assign mem[4025] = 5'h02;
  assign mem[4026] = 5'h11;
  assign mem[4027] = 5'h10;
  assign mem[4028] = 5'h00;
  assign mem[4029] = 5'h01;
  assign mem[4030] = 5'h10;
  assign mem[4031] = 5'h00;
  assign mem[4032] = 5'h05;
  assign mem[4033] = 5'h14;
  assign mem[4034] = 5'h13;
  assign mem[4035] = 5'h12;
  assign mem[4036] = 5'h11;
  assign mem[4037] = 5'h10;
  assign mem[4038] = 5'h00;
  assign mem[4039] = 5'h01;
  assign mem[4040] = 5'h10;
  assign mem[4041] = 5'h00;
  assign mem[4042] = 5'h02;
  assign mem[4043] = 5'h11;
  assign mem[4044] = 5'h10;
  assign mem[4045] = 5'h00;
  assign mem[4046] = 5'h01;
  assign mem[4047] = 5'h10;
  assign mem[4048] = 5'h00;
  assign mem[4049] = 5'h03;
  assign mem[4050] = 5'h12;
  assign mem[4051] = 5'h11;
  assign mem[4052] = 5'h10;
  assign mem[4053] = 5'h00;
  assign mem[4054] = 5'h01;
  assign mem[4055] = 5'h10;
  assign mem[4056] = 5'h00;
  assign mem[4057] = 5'h02;
  assign mem[4058] = 5'h11;
  assign mem[4059] = 5'h10;
  assign mem[4060] = 5'h00;
  assign mem[4061] = 5'h01;
  assign mem[4062] = 5'h10;
  assign mem[4063] = 5'h00;
  assign mem[4064] = 5'h04;
  assign mem[4065] = 5'h13;
  assign mem[4066] = 5'h12;
  assign mem[4067] = 5'h11;
  assign mem[4068] = 5'h10;
  assign mem[4069] = 5'h00;
  assign mem[4070] = 5'h01;
  assign mem[4071] = 5'h10;
  assign mem[4072] = 5'h00;
  assign mem[4073] = 5'h02;
  assign mem[4074] = 5'h11;
  assign mem[4075] = 5'h10;
  assign mem[4076] = 5'h00;
  assign mem[4077] = 5'h01;
  assign mem[4078] = 5'h10;
  assign mem[4079] = 5'h00;
  assign mem[4080] = 5'h03;
  assign mem[4081] = 5'h12;
  assign mem[4082] = 5'h11;
  assign mem[4083] = 5'h10;
  assign mem[4084] = 5'h00;
  assign mem[4085] = 5'h01;
  assign mem[4086] = 5'h10;
  assign mem[4087] = 5'h00;
  assign mem[4088] = 5'h02;
  assign mem[4089] = 5'h11;
  assign mem[4090] = 5'h10;
  assign mem[4091] = 5'h00;
  assign mem[4092] = 5'h01;
  assign mem[4093] = 5'h10;
  assign mem[4094] = 5'h00;
  assign mem[4095] = 5'h0b;
  assign mem[4096] = 5'h1a;
  assign mem[4097] = 5'h19;
  assign mem[4098] = 5'h18;
  assign mem[4099] = 5'h17;
  assign mem[4100] = 5'h16;
  assign mem[4101] = 5'h15;
  assign mem[4102] = 5'h14;
  assign mem[4103] = 5'h13;
  assign mem[4104] = 5'h12;
  assign mem[4105] = 5'h11;
  assign mem[4106] = 5'h10;
  assign mem[4107] = 5'h00;
  assign mem[4108] = 5'h01;
  assign mem[4109] = 5'h10;
  assign mem[4110] = 5'h00;
  assign mem[4111] = 5'h02;
  assign mem[4112] = 5'h11;
  assign mem[4113] = 5'h10;
  assign mem[4114] = 5'h00;
  assign mem[4115] = 5'h01;
  assign mem[4116] = 5'h10;
  assign mem[4117] = 5'h00;
  assign mem[4118] = 5'h03;
  assign mem[4119] = 5'h12;
  assign mem[4120] = 5'h11;
  assign mem[4121] = 5'h10;
  assign mem[4122] = 5'h00;
  assign mem[4123] = 5'h01;
  assign mem[4124] = 5'h10;
  assign mem[4125] = 5'h00;
  assign mem[4126] = 5'h02;
  assign mem[4127] = 5'h11;
  assign mem[4128] = 5'h10;
  assign mem[4129] = 5'h00;
  assign mem[4130] = 5'h01;
  assign mem[4131] = 5'h10;
  assign mem[4132] = 5'h00;
  assign mem[4133] = 5'h04;
  assign mem[4134] = 5'h13;
  assign mem[4135] = 5'h12;
  assign mem[4136] = 5'h11;
  assign mem[4137] = 5'h10;
  assign mem[4138] = 5'h00;
  assign mem[4139] = 5'h01;
  assign mem[4140] = 5'h10;
  assign mem[4141] = 5'h00;
  assign mem[4142] = 5'h02;
  assign mem[4143] = 5'h11;
  assign mem[4144] = 5'h10;
  assign mem[4145] = 5'h00;
  assign mem[4146] = 5'h01;
  assign mem[4147] = 5'h10;
  assign mem[4148] = 5'h00;
  assign mem[4149] = 5'h03;
  assign mem[4150] = 5'h12;
  assign mem[4151] = 5'h11;
  assign mem[4152] = 5'h10;
  assign mem[4153] = 5'h00;
  assign mem[4154] = 5'h01;
  assign mem[4155] = 5'h10;
  assign mem[4156] = 5'h00;
  assign mem[4157] = 5'h02;
  assign mem[4158] = 5'h11;
  assign mem[4159] = 5'h10;
  assign mem[4160] = 5'h00;
  assign mem[4161] = 5'h01;
  assign mem[4162] = 5'h10;
  assign mem[4163] = 5'h00;
  assign mem[4164] = 5'h05;
  assign mem[4165] = 5'h14;
  assign mem[4166] = 5'h13;
  assign mem[4167] = 5'h12;
  assign mem[4168] = 5'h11;
  assign mem[4169] = 5'h10;
  assign mem[4170] = 5'h00;
  assign mem[4171] = 5'h01;
  assign mem[4172] = 5'h10;
  assign mem[4173] = 5'h00;
  assign mem[4174] = 5'h02;
  assign mem[4175] = 5'h11;
  assign mem[4176] = 5'h10;
  assign mem[4177] = 5'h00;
  assign mem[4178] = 5'h01;
  assign mem[4179] = 5'h10;
  assign mem[4180] = 5'h00;
  assign mem[4181] = 5'h03;
  assign mem[4182] = 5'h12;
  assign mem[4183] = 5'h11;
  assign mem[4184] = 5'h10;
  assign mem[4185] = 5'h00;
  assign mem[4186] = 5'h01;
  assign mem[4187] = 5'h10;
  assign mem[4188] = 5'h00;
  assign mem[4189] = 5'h02;
  assign mem[4190] = 5'h11;
  assign mem[4191] = 5'h10;
  assign mem[4192] = 5'h00;
  assign mem[4193] = 5'h01;
  assign mem[4194] = 5'h10;
  assign mem[4195] = 5'h00;
  assign mem[4196] = 5'h04;
  assign mem[4197] = 5'h13;
  assign mem[4198] = 5'h12;
  assign mem[4199] = 5'h11;
  assign mem[4200] = 5'h10;
  assign mem[4201] = 5'h00;
  assign mem[4202] = 5'h01;
  assign mem[4203] = 5'h10;
  assign mem[4204] = 5'h00;
  assign mem[4205] = 5'h02;
  assign mem[4206] = 5'h11;
  assign mem[4207] = 5'h10;
  assign mem[4208] = 5'h00;
  assign mem[4209] = 5'h01;
  assign mem[4210] = 5'h10;
  assign mem[4211] = 5'h00;
  assign mem[4212] = 5'h03;
  assign mem[4213] = 5'h12;
  assign mem[4214] = 5'h11;
  assign mem[4215] = 5'h10;
  assign mem[4216] = 5'h00;
  assign mem[4217] = 5'h01;
  assign mem[4218] = 5'h10;
  assign mem[4219] = 5'h00;
  assign mem[4220] = 5'h02;
  assign mem[4221] = 5'h11;
  assign mem[4222] = 5'h10;
  assign mem[4223] = 5'h00;
  assign mem[4224] = 5'h01;
  assign mem[4225] = 5'h10;
  assign mem[4226] = 5'h00;
  assign mem[4227] = 5'h06;
  assign mem[4228] = 5'h15;
  assign mem[4229] = 5'h14;
  assign mem[4230] = 5'h13;
  assign mem[4231] = 5'h12;
  assign mem[4232] = 5'h11;
  assign mem[4233] = 5'h10;
  assign mem[4234] = 5'h00;
  assign mem[4235] = 5'h01;
  assign mem[4236] = 5'h10;
  assign mem[4237] = 5'h00;
  assign mem[4238] = 5'h02;
  assign mem[4239] = 5'h11;
  assign mem[4240] = 5'h10;
  assign mem[4241] = 5'h00;
  assign mem[4242] = 5'h01;
  assign mem[4243] = 5'h10;
  assign mem[4244] = 5'h00;
  assign mem[4245] = 5'h03;
  assign mem[4246] = 5'h12;
  assign mem[4247] = 5'h11;
  assign mem[4248] = 5'h10;
  assign mem[4249] = 5'h00;
  assign mem[4250] = 5'h01;
  assign mem[4251] = 5'h10;
  assign mem[4252] = 5'h00;
  assign mem[4253] = 5'h02;
  assign mem[4254] = 5'h11;
  assign mem[4255] = 5'h10;
  assign mem[4256] = 5'h00;
  assign mem[4257] = 5'h01;
  assign mem[4258] = 5'h10;
  assign mem[4259] = 5'h00;
  assign mem[4260] = 5'h04;
  assign mem[4261] = 5'h13;
  assign mem[4262] = 5'h12;
  assign mem[4263] = 5'h11;
  assign mem[4264] = 5'h10;
  assign mem[4265] = 5'h00;
  assign mem[4266] = 5'h01;
  assign mem[4267] = 5'h10;
  assign mem[4268] = 5'h00;
  assign mem[4269] = 5'h02;
  assign mem[4270] = 5'h11;
  assign mem[4271] = 5'h10;
  assign mem[4272] = 5'h00;
  assign mem[4273] = 5'h01;
  assign mem[4274] = 5'h10;
  assign mem[4275] = 5'h00;
  assign mem[4276] = 5'h03;
  assign mem[4277] = 5'h12;
  assign mem[4278] = 5'h11;
  assign mem[4279] = 5'h10;
  assign mem[4280] = 5'h00;
  assign mem[4281] = 5'h01;
  assign mem[4282] = 5'h10;
  assign mem[4283] = 5'h00;
  assign mem[4284] = 5'h02;
  assign mem[4285] = 5'h11;
  assign mem[4286] = 5'h10;
  assign mem[4287] = 5'h00;
  assign mem[4288] = 5'h01;
  assign mem[4289] = 5'h10;
  assign mem[4290] = 5'h00;
  assign mem[4291] = 5'h05;
  assign mem[4292] = 5'h14;
  assign mem[4293] = 5'h13;
  assign mem[4294] = 5'h12;
  assign mem[4295] = 5'h11;
  assign mem[4296] = 5'h10;
  assign mem[4297] = 5'h00;
  assign mem[4298] = 5'h01;
  assign mem[4299] = 5'h10;
  assign mem[4300] = 5'h00;
  assign mem[4301] = 5'h02;
  assign mem[4302] = 5'h11;
  assign mem[4303] = 5'h10;
  assign mem[4304] = 5'h00;
  assign mem[4305] = 5'h01;
  assign mem[4306] = 5'h10;
  assign mem[4307] = 5'h00;
  assign mem[4308] = 5'h03;
  assign mem[4309] = 5'h12;
  assign mem[4310] = 5'h11;
  assign mem[4311] = 5'h10;
  assign mem[4312] = 5'h00;
  assign mem[4313] = 5'h01;
  assign mem[4314] = 5'h10;
  assign mem[4315] = 5'h00;
  assign mem[4316] = 5'h02;
  assign mem[4317] = 5'h11;
  assign mem[4318] = 5'h10;
  assign mem[4319] = 5'h00;
  assign mem[4320] = 5'h01;
  assign mem[4321] = 5'h10;
  assign mem[4322] = 5'h00;
  assign mem[4323] = 5'h04;
  assign mem[4324] = 5'h13;
  assign mem[4325] = 5'h12;
  assign mem[4326] = 5'h11;
  assign mem[4327] = 5'h10;
  assign mem[4328] = 5'h00;
  assign mem[4329] = 5'h01;
  assign mem[4330] = 5'h10;
  assign mem[4331] = 5'h00;
  assign mem[4332] = 5'h02;
  assign mem[4333] = 5'h11;
  assign mem[4334] = 5'h10;
  assign mem[4335] = 5'h00;
  assign mem[4336] = 5'h01;
  assign mem[4337] = 5'h10;
  assign mem[4338] = 5'h00;
  assign mem[4339] = 5'h03;
  assign mem[4340] = 5'h12;
  assign mem[4341] = 5'h11;
  assign mem[4342] = 5'h10;
  assign mem[4343] = 5'h00;
  assign mem[4344] = 5'h01;
  assign mem[4345] = 5'h10;
  assign mem[4346] = 5'h00;
  assign mem[4347] = 5'h02;
  assign mem[4348] = 5'h11;
  assign mem[4349] = 5'h10;
  assign mem[4350] = 5'h00;
  assign mem[4351] = 5'h01;
  assign mem[4352] = 5'h10;
  assign mem[4353] = 5'h00;
  assign mem[4354] = 5'h07;
  assign mem[4355] = 5'h16;
  assign mem[4356] = 5'h15;
  assign mem[4357] = 5'h14;
  assign mem[4358] = 5'h13;
  assign mem[4359] = 5'h12;
  assign mem[4360] = 5'h11;
  assign mem[4361] = 5'h10;
  assign mem[4362] = 5'h00;
  assign mem[4363] = 5'h01;
  assign mem[4364] = 5'h10;
  assign mem[4365] = 5'h00;
  assign mem[4366] = 5'h02;
  assign mem[4367] = 5'h11;
  assign mem[4368] = 5'h10;
  assign mem[4369] = 5'h00;
  assign mem[4370] = 5'h01;
  assign mem[4371] = 5'h10;
  assign mem[4372] = 5'h00;
  assign mem[4373] = 5'h03;
  assign mem[4374] = 5'h12;
  assign mem[4375] = 5'h11;
  assign mem[4376] = 5'h10;
  assign mem[4377] = 5'h00;
  assign mem[4378] = 5'h01;
  assign mem[4379] = 5'h10;
  assign mem[4380] = 5'h00;
  assign mem[4381] = 5'h02;
  assign mem[4382] = 5'h11;
  assign mem[4383] = 5'h10;
  assign mem[4384] = 5'h00;
  assign mem[4385] = 5'h01;
  assign mem[4386] = 5'h10;
  assign mem[4387] = 5'h00;
  assign mem[4388] = 5'h04;
  assign mem[4389] = 5'h13;
  assign mem[4390] = 5'h12;
  assign mem[4391] = 5'h11;
  assign mem[4392] = 5'h10;
  assign mem[4393] = 5'h00;
  assign mem[4394] = 5'h01;
  assign mem[4395] = 5'h10;
  assign mem[4396] = 5'h00;
  assign mem[4397] = 5'h02;
  assign mem[4398] = 5'h11;
  assign mem[4399] = 5'h10;
  assign mem[4400] = 5'h00;
  assign mem[4401] = 5'h01;
  assign mem[4402] = 5'h10;
  assign mem[4403] = 5'h00;
  assign mem[4404] = 5'h03;
  assign mem[4405] = 5'h12;
  assign mem[4406] = 5'h11;
  assign mem[4407] = 5'h10;
  assign mem[4408] = 5'h00;
  assign mem[4409] = 5'h01;
  assign mem[4410] = 5'h10;
  assign mem[4411] = 5'h00;
  assign mem[4412] = 5'h02;
  assign mem[4413] = 5'h11;
  assign mem[4414] = 5'h10;
  assign mem[4415] = 5'h00;
  assign mem[4416] = 5'h01;
  assign mem[4417] = 5'h10;
  assign mem[4418] = 5'h00;
  assign mem[4419] = 5'h05;
  assign mem[4420] = 5'h14;
  assign mem[4421] = 5'h13;
  assign mem[4422] = 5'h12;
  assign mem[4423] = 5'h11;
  assign mem[4424] = 5'h10;
  assign mem[4425] = 5'h00;
  assign mem[4426] = 5'h01;
  assign mem[4427] = 5'h10;
  assign mem[4428] = 5'h00;
  assign mem[4429] = 5'h02;
  assign mem[4430] = 5'h11;
  assign mem[4431] = 5'h10;
  assign mem[4432] = 5'h00;
  assign mem[4433] = 5'h01;
  assign mem[4434] = 5'h10;
  assign mem[4435] = 5'h00;
  assign mem[4436] = 5'h03;
  assign mem[4437] = 5'h12;
  assign mem[4438] = 5'h11;
  assign mem[4439] = 5'h10;
  assign mem[4440] = 5'h00;
  assign mem[4441] = 5'h01;
  assign mem[4442] = 5'h10;
  assign mem[4443] = 5'h00;
  assign mem[4444] = 5'h02;
  assign mem[4445] = 5'h11;
  assign mem[4446] = 5'h10;
  assign mem[4447] = 5'h00;
  assign mem[4448] = 5'h01;
  assign mem[4449] = 5'h10;
  assign mem[4450] = 5'h00;
  assign mem[4451] = 5'h04;
  assign mem[4452] = 5'h13;
  assign mem[4453] = 5'h12;
  assign mem[4454] = 5'h11;
  assign mem[4455] = 5'h10;
  assign mem[4456] = 5'h00;
  assign mem[4457] = 5'h01;
  assign mem[4458] = 5'h10;
  assign mem[4459] = 5'h00;
  assign mem[4460] = 5'h02;
  assign mem[4461] = 5'h11;
  assign mem[4462] = 5'h10;
  assign mem[4463] = 5'h00;
  assign mem[4464] = 5'h01;
  assign mem[4465] = 5'h10;
  assign mem[4466] = 5'h00;
  assign mem[4467] = 5'h03;
  assign mem[4468] = 5'h12;
  assign mem[4469] = 5'h11;
  assign mem[4470] = 5'h10;
  assign mem[4471] = 5'h00;
  assign mem[4472] = 5'h01;
  assign mem[4473] = 5'h10;
  assign mem[4474] = 5'h00;
  assign mem[4475] = 5'h02;
  assign mem[4476] = 5'h11;
  assign mem[4477] = 5'h10;
  assign mem[4478] = 5'h00;
  assign mem[4479] = 5'h01;
  assign mem[4480] = 5'h10;
  assign mem[4481] = 5'h00;
  assign mem[4482] = 5'h06;
  assign mem[4483] = 5'h15;
  assign mem[4484] = 5'h14;
  assign mem[4485] = 5'h13;
  assign mem[4486] = 5'h12;
  assign mem[4487] = 5'h11;
  assign mem[4488] = 5'h10;
  assign mem[4489] = 5'h00;
  assign mem[4490] = 5'h01;
  assign mem[4491] = 5'h10;
  assign mem[4492] = 5'h00;
  assign mem[4493] = 5'h02;
  assign mem[4494] = 5'h11;
  assign mem[4495] = 5'h10;
  assign mem[4496] = 5'h00;
  assign mem[4497] = 5'h01;
  assign mem[4498] = 5'h10;
  assign mem[4499] = 5'h00;
  assign mem[4500] = 5'h03;
  assign mem[4501] = 5'h12;
  assign mem[4502] = 5'h11;
  assign mem[4503] = 5'h10;
  assign mem[4504] = 5'h00;
  assign mem[4505] = 5'h01;
  assign mem[4506] = 5'h10;
  assign mem[4507] = 5'h00;
  assign mem[4508] = 5'h02;
  assign mem[4509] = 5'h11;
  assign mem[4510] = 5'h10;
  assign mem[4511] = 5'h00;
  assign mem[4512] = 5'h01;
  assign mem[4513] = 5'h10;
  assign mem[4514] = 5'h00;
  assign mem[4515] = 5'h04;
  assign mem[4516] = 5'h13;
  assign mem[4517] = 5'h12;
  assign mem[4518] = 5'h11;
  assign mem[4519] = 5'h10;
  assign mem[4520] = 5'h00;
  assign mem[4521] = 5'h01;
  assign mem[4522] = 5'h10;
  assign mem[4523] = 5'h00;
  assign mem[4524] = 5'h02;
  assign mem[4525] = 5'h11;
  assign mem[4526] = 5'h10;
  assign mem[4527] = 5'h00;
  assign mem[4528] = 5'h01;
  assign mem[4529] = 5'h10;
  assign mem[4530] = 5'h00;
  assign mem[4531] = 5'h03;
  assign mem[4532] = 5'h12;
  assign mem[4533] = 5'h11;
  assign mem[4534] = 5'h10;
  assign mem[4535] = 5'h00;
  assign mem[4536] = 5'h01;
  assign mem[4537] = 5'h10;
  assign mem[4538] = 5'h00;
  assign mem[4539] = 5'h02;
  assign mem[4540] = 5'h11;
  assign mem[4541] = 5'h10;
  assign mem[4542] = 5'h00;
  assign mem[4543] = 5'h01;
  assign mem[4544] = 5'h10;
  assign mem[4545] = 5'h00;
  assign mem[4546] = 5'h05;
  assign mem[4547] = 5'h14;
  assign mem[4548] = 5'h13;
  assign mem[4549] = 5'h12;
  assign mem[4550] = 5'h11;
  assign mem[4551] = 5'h10;
  assign mem[4552] = 5'h00;
  assign mem[4553] = 5'h01;
  assign mem[4554] = 5'h10;
  assign mem[4555] = 5'h00;
  assign mem[4556] = 5'h02;
  assign mem[4557] = 5'h11;
  assign mem[4558] = 5'h10;
  assign mem[4559] = 5'h00;
  assign mem[4560] = 5'h01;
  assign mem[4561] = 5'h10;
  assign mem[4562] = 5'h00;
  assign mem[4563] = 5'h03;
  assign mem[4564] = 5'h12;
  assign mem[4565] = 5'h11;
  assign mem[4566] = 5'h10;
  assign mem[4567] = 5'h00;
  assign mem[4568] = 5'h01;
  assign mem[4569] = 5'h10;
  assign mem[4570] = 5'h00;
  assign mem[4571] = 5'h02;
  assign mem[4572] = 5'h11;
  assign mem[4573] = 5'h10;
  assign mem[4574] = 5'h00;
  assign mem[4575] = 5'h01;
  assign mem[4576] = 5'h10;
  assign mem[4577] = 5'h00;
  assign mem[4578] = 5'h04;
  assign mem[4579] = 5'h13;
  assign mem[4580] = 5'h12;
  assign mem[4581] = 5'h11;
  assign mem[4582] = 5'h10;
  assign mem[4583] = 5'h00;
  assign mem[4584] = 5'h01;
  assign mem[4585] = 5'h10;
  assign mem[4586] = 5'h00;
  assign mem[4587] = 5'h02;
  assign mem[4588] = 5'h11;
  assign mem[4589] = 5'h10;
  assign mem[4590] = 5'h00;
  assign mem[4591] = 5'h01;
  assign mem[4592] = 5'h10;
  assign mem[4593] = 5'h00;
  assign mem[4594] = 5'h03;
  assign mem[4595] = 5'h12;
  assign mem[4596] = 5'h11;
  assign mem[4597] = 5'h10;
  assign mem[4598] = 5'h00;
  assign mem[4599] = 5'h01;
  assign mem[4600] = 5'h10;
  assign mem[4601] = 5'h00;
  assign mem[4602] = 5'h02;
  assign mem[4603] = 5'h11;
  assign mem[4604] = 5'h10;
  assign mem[4605] = 5'h00;
  assign mem[4606] = 5'h01;
  assign mem[4607] = 5'h10;
  assign mem[4608] = 5'h00;
  assign mem[4609] = 5'h08;
  assign mem[4610] = 5'h17;
  assign mem[4611] = 5'h16;
  assign mem[4612] = 5'h15;
  assign mem[4613] = 5'h14;
  assign mem[4614] = 5'h13;
  assign mem[4615] = 5'h12;
  assign mem[4616] = 5'h11;
  assign mem[4617] = 5'h10;
  assign mem[4618] = 5'h00;
  assign mem[4619] = 5'h01;
  assign mem[4620] = 5'h10;
  assign mem[4621] = 5'h00;
  assign mem[4622] = 5'h02;
  assign mem[4623] = 5'h11;
  assign mem[4624] = 5'h10;
  assign mem[4625] = 5'h00;
  assign mem[4626] = 5'h01;
  assign mem[4627] = 5'h10;
  assign mem[4628] = 5'h00;
  assign mem[4629] = 5'h03;
  assign mem[4630] = 5'h12;
  assign mem[4631] = 5'h11;
  assign mem[4632] = 5'h10;
  assign mem[4633] = 5'h00;
  assign mem[4634] = 5'h01;
  assign mem[4635] = 5'h10;
  assign mem[4636] = 5'h00;
  assign mem[4637] = 5'h02;
  assign mem[4638] = 5'h11;
  assign mem[4639] = 5'h10;
  assign mem[4640] = 5'h00;
  assign mem[4641] = 5'h01;
  assign mem[4642] = 5'h10;
  assign mem[4643] = 5'h00;
  assign mem[4644] = 5'h04;
  assign mem[4645] = 5'h13;
  assign mem[4646] = 5'h12;
  assign mem[4647] = 5'h11;
  assign mem[4648] = 5'h10;
  assign mem[4649] = 5'h00;
  assign mem[4650] = 5'h01;
  assign mem[4651] = 5'h10;
  assign mem[4652] = 5'h00;
  assign mem[4653] = 5'h02;
  assign mem[4654] = 5'h11;
  assign mem[4655] = 5'h10;
  assign mem[4656] = 5'h00;
  assign mem[4657] = 5'h01;
  assign mem[4658] = 5'h10;
  assign mem[4659] = 5'h00;
  assign mem[4660] = 5'h03;
  assign mem[4661] = 5'h12;
  assign mem[4662] = 5'h11;
  assign mem[4663] = 5'h10;
  assign mem[4664] = 5'h00;
  assign mem[4665] = 5'h01;
  assign mem[4666] = 5'h10;
  assign mem[4667] = 5'h00;
  assign mem[4668] = 5'h02;
  assign mem[4669] = 5'h11;
  assign mem[4670] = 5'h10;
  assign mem[4671] = 5'h00;
  assign mem[4672] = 5'h01;
  assign mem[4673] = 5'h10;
  assign mem[4674] = 5'h00;
  assign mem[4675] = 5'h05;
  assign mem[4676] = 5'h14;
  assign mem[4677] = 5'h13;
  assign mem[4678] = 5'h12;
  assign mem[4679] = 5'h11;
  assign mem[4680] = 5'h10;
  assign mem[4681] = 5'h00;
  assign mem[4682] = 5'h01;
  assign mem[4683] = 5'h10;
  assign mem[4684] = 5'h00;
  assign mem[4685] = 5'h02;
  assign mem[4686] = 5'h11;
  assign mem[4687] = 5'h10;
  assign mem[4688] = 5'h00;
  assign mem[4689] = 5'h01;
  assign mem[4690] = 5'h10;
  assign mem[4691] = 5'h00;
  assign mem[4692] = 5'h03;
  assign mem[4693] = 5'h12;
  assign mem[4694] = 5'h11;
  assign mem[4695] = 5'h10;
  assign mem[4696] = 5'h00;
  assign mem[4697] = 5'h01;
  assign mem[4698] = 5'h10;
  assign mem[4699] = 5'h00;
  assign mem[4700] = 5'h02;
  assign mem[4701] = 5'h11;
  assign mem[4702] = 5'h10;
  assign mem[4703] = 5'h00;
  assign mem[4704] = 5'h01;
  assign mem[4705] = 5'h10;
  assign mem[4706] = 5'h00;
  assign mem[4707] = 5'h04;
  assign mem[4708] = 5'h13;
  assign mem[4709] = 5'h12;
  assign mem[4710] = 5'h11;
  assign mem[4711] = 5'h10;
  assign mem[4712] = 5'h00;
  assign mem[4713] = 5'h01;
  assign mem[4714] = 5'h10;
  assign mem[4715] = 5'h00;
  assign mem[4716] = 5'h02;
  assign mem[4717] = 5'h11;
  assign mem[4718] = 5'h10;
  assign mem[4719] = 5'h00;
  assign mem[4720] = 5'h01;
  assign mem[4721] = 5'h10;
  assign mem[4722] = 5'h00;
  assign mem[4723] = 5'h03;
  assign mem[4724] = 5'h12;
  assign mem[4725] = 5'h11;
  assign mem[4726] = 5'h10;
  assign mem[4727] = 5'h00;
  assign mem[4728] = 5'h01;
  assign mem[4729] = 5'h10;
  assign mem[4730] = 5'h00;
  assign mem[4731] = 5'h02;
  assign mem[4732] = 5'h11;
  assign mem[4733] = 5'h10;
  assign mem[4734] = 5'h00;
  assign mem[4735] = 5'h01;
  assign mem[4736] = 5'h10;
  assign mem[4737] = 5'h00;
  assign mem[4738] = 5'h06;
  assign mem[4739] = 5'h15;
  assign mem[4740] = 5'h14;
  assign mem[4741] = 5'h13;
  assign mem[4742] = 5'h12;
  assign mem[4743] = 5'h11;
  assign mem[4744] = 5'h10;
  assign mem[4745] = 5'h00;
  assign mem[4746] = 5'h01;
  assign mem[4747] = 5'h10;
  assign mem[4748] = 5'h00;
  assign mem[4749] = 5'h02;
  assign mem[4750] = 5'h11;
  assign mem[4751] = 5'h10;
  assign mem[4752] = 5'h00;
  assign mem[4753] = 5'h01;
  assign mem[4754] = 5'h10;
  assign mem[4755] = 5'h00;
  assign mem[4756] = 5'h03;
  assign mem[4757] = 5'h12;
  assign mem[4758] = 5'h11;
  assign mem[4759] = 5'h10;
  assign mem[4760] = 5'h00;
  assign mem[4761] = 5'h01;
  assign mem[4762] = 5'h10;
  assign mem[4763] = 5'h00;
  assign mem[4764] = 5'h02;
  assign mem[4765] = 5'h11;
  assign mem[4766] = 5'h10;
  assign mem[4767] = 5'h00;
  assign mem[4768] = 5'h01;
  assign mem[4769] = 5'h10;
  assign mem[4770] = 5'h00;
  assign mem[4771] = 5'h04;
  assign mem[4772] = 5'h13;
  assign mem[4773] = 5'h12;
  assign mem[4774] = 5'h11;
  assign mem[4775] = 5'h10;
  assign mem[4776] = 5'h00;
  assign mem[4777] = 5'h01;
  assign mem[4778] = 5'h10;
  assign mem[4779] = 5'h00;
  assign mem[4780] = 5'h02;
  assign mem[4781] = 5'h11;
  assign mem[4782] = 5'h10;
  assign mem[4783] = 5'h00;
  assign mem[4784] = 5'h01;
  assign mem[4785] = 5'h10;
  assign mem[4786] = 5'h00;
  assign mem[4787] = 5'h03;
  assign mem[4788] = 5'h12;
  assign mem[4789] = 5'h11;
  assign mem[4790] = 5'h10;
  assign mem[4791] = 5'h00;
  assign mem[4792] = 5'h01;
  assign mem[4793] = 5'h10;
  assign mem[4794] = 5'h00;
  assign mem[4795] = 5'h02;
  assign mem[4796] = 5'h11;
  assign mem[4797] = 5'h10;
  assign mem[4798] = 5'h00;
  assign mem[4799] = 5'h01;
  assign mem[4800] = 5'h10;
  assign mem[4801] = 5'h00;
  assign mem[4802] = 5'h05;
  assign mem[4803] = 5'h14;
  assign mem[4804] = 5'h13;
  assign mem[4805] = 5'h12;
  assign mem[4806] = 5'h11;
  assign mem[4807] = 5'h10;
  assign mem[4808] = 5'h00;
  assign mem[4809] = 5'h01;
  assign mem[4810] = 5'h10;
  assign mem[4811] = 5'h00;
  assign mem[4812] = 5'h02;
  assign mem[4813] = 5'h11;
  assign mem[4814] = 5'h10;
  assign mem[4815] = 5'h00;
  assign mem[4816] = 5'h01;
  assign mem[4817] = 5'h10;
  assign mem[4818] = 5'h00;
  assign mem[4819] = 5'h03;
  assign mem[4820] = 5'h12;
  assign mem[4821] = 5'h11;
  assign mem[4822] = 5'h10;
  assign mem[4823] = 5'h00;
  assign mem[4824] = 5'h01;
  assign mem[4825] = 5'h10;
  assign mem[4826] = 5'h00;
  assign mem[4827] = 5'h02;
  assign mem[4828] = 5'h11;
  assign mem[4829] = 5'h10;
  assign mem[4830] = 5'h00;
  assign mem[4831] = 5'h01;
  assign mem[4832] = 5'h10;
  assign mem[4833] = 5'h00;
  assign mem[4834] = 5'h04;
  assign mem[4835] = 5'h13;
  assign mem[4836] = 5'h12;
  assign mem[4837] = 5'h11;
  assign mem[4838] = 5'h10;
  assign mem[4839] = 5'h00;
  assign mem[4840] = 5'h01;
  assign mem[4841] = 5'h10;
  assign mem[4842] = 5'h00;
  assign mem[4843] = 5'h02;
  assign mem[4844] = 5'h11;
  assign mem[4845] = 5'h10;
  assign mem[4846] = 5'h00;
  assign mem[4847] = 5'h01;
  assign mem[4848] = 5'h10;
  assign mem[4849] = 5'h00;
  assign mem[4850] = 5'h03;
  assign mem[4851] = 5'h12;
  assign mem[4852] = 5'h11;
  assign mem[4853] = 5'h10;
  assign mem[4854] = 5'h00;
  assign mem[4855] = 5'h01;
  assign mem[4856] = 5'h10;
  assign mem[4857] = 5'h00;
  assign mem[4858] = 5'h02;
  assign mem[4859] = 5'h11;
  assign mem[4860] = 5'h10;
  assign mem[4861] = 5'h00;
  assign mem[4862] = 5'h01;
  assign mem[4863] = 5'h10;
  assign mem[4864] = 5'h00;
  assign mem[4865] = 5'h07;
  assign mem[4866] = 5'h16;
  assign mem[4867] = 5'h15;
  assign mem[4868] = 5'h14;
  assign mem[4869] = 5'h13;
  assign mem[4870] = 5'h12;
  assign mem[4871] = 5'h11;
  assign mem[4872] = 5'h10;
  assign mem[4873] = 5'h00;
  assign mem[4874] = 5'h01;
  assign mem[4875] = 5'h10;
  assign mem[4876] = 5'h00;
  assign mem[4877] = 5'h02;
  assign mem[4878] = 5'h11;
  assign mem[4879] = 5'h10;
  assign mem[4880] = 5'h00;
  assign mem[4881] = 5'h01;
  assign mem[4882] = 5'h10;
  assign mem[4883] = 5'h00;
  assign mem[4884] = 5'h03;
  assign mem[4885] = 5'h12;
  assign mem[4886] = 5'h11;
  assign mem[4887] = 5'h10;
  assign mem[4888] = 5'h00;
  assign mem[4889] = 5'h01;
  assign mem[4890] = 5'h10;
  assign mem[4891] = 5'h00;
  assign mem[4892] = 5'h02;
  assign mem[4893] = 5'h11;
  assign mem[4894] = 5'h10;
  assign mem[4895] = 5'h00;
  assign mem[4896] = 5'h01;
  assign mem[4897] = 5'h10;
  assign mem[4898] = 5'h00;
  assign mem[4899] = 5'h04;
  assign mem[4900] = 5'h13;
  assign mem[4901] = 5'h12;
  assign mem[4902] = 5'h11;
  assign mem[4903] = 5'h10;
  assign mem[4904] = 5'h00;
  assign mem[4905] = 5'h01;
  assign mem[4906] = 5'h10;
  assign mem[4907] = 5'h00;
  assign mem[4908] = 5'h02;
  assign mem[4909] = 5'h11;
  assign mem[4910] = 5'h10;
  assign mem[4911] = 5'h00;
  assign mem[4912] = 5'h01;
  assign mem[4913] = 5'h10;
  assign mem[4914] = 5'h00;
  assign mem[4915] = 5'h03;
  assign mem[4916] = 5'h12;
  assign mem[4917] = 5'h11;
  assign mem[4918] = 5'h10;
  assign mem[4919] = 5'h00;
  assign mem[4920] = 5'h01;
  assign mem[4921] = 5'h10;
  assign mem[4922] = 5'h00;
  assign mem[4923] = 5'h02;
  assign mem[4924] = 5'h11;
  assign mem[4925] = 5'h10;
  assign mem[4926] = 5'h00;
  assign mem[4927] = 5'h01;
  assign mem[4928] = 5'h10;
  assign mem[4929] = 5'h00;
  assign mem[4930] = 5'h05;
  assign mem[4931] = 5'h14;
  assign mem[4932] = 5'h13;
  assign mem[4933] = 5'h12;
  assign mem[4934] = 5'h11;
  assign mem[4935] = 5'h10;
  assign mem[4936] = 5'h00;
  assign mem[4937] = 5'h01;
  assign mem[4938] = 5'h10;
  assign mem[4939] = 5'h00;
  assign mem[4940] = 5'h02;
  assign mem[4941] = 5'h11;
  assign mem[4942] = 5'h10;
  assign mem[4943] = 5'h00;
  assign mem[4944] = 5'h01;
  assign mem[4945] = 5'h10;
  assign mem[4946] = 5'h00;
  assign mem[4947] = 5'h03;
  assign mem[4948] = 5'h12;
  assign mem[4949] = 5'h11;
  assign mem[4950] = 5'h10;
  assign mem[4951] = 5'h00;
  assign mem[4952] = 5'h01;
  assign mem[4953] = 5'h10;
  assign mem[4954] = 5'h00;
  assign mem[4955] = 5'h02;
  assign mem[4956] = 5'h11;
  assign mem[4957] = 5'h10;
  assign mem[4958] = 5'h00;
  assign mem[4959] = 5'h01;
  assign mem[4960] = 5'h10;
  assign mem[4961] = 5'h00;
  assign mem[4962] = 5'h04;
  assign mem[4963] = 5'h13;
  assign mem[4964] = 5'h12;
  assign mem[4965] = 5'h11;
  assign mem[4966] = 5'h10;
  assign mem[4967] = 5'h00;
  assign mem[4968] = 5'h01;
  assign mem[4969] = 5'h10;
  assign mem[4970] = 5'h00;
  assign mem[4971] = 5'h02;
  assign mem[4972] = 5'h11;
  assign mem[4973] = 5'h10;
  assign mem[4974] = 5'h00;
  assign mem[4975] = 5'h01;
  assign mem[4976] = 5'h10;
  assign mem[4977] = 5'h00;
  assign mem[4978] = 5'h03;
  assign mem[4979] = 5'h12;
  assign mem[4980] = 5'h11;
  assign mem[4981] = 5'h10;
  assign mem[4982] = 5'h00;
  assign mem[4983] = 5'h01;
  assign mem[4984] = 5'h10;
  assign mem[4985] = 5'h00;
  assign mem[4986] = 5'h02;
  assign mem[4987] = 5'h11;
  assign mem[4988] = 5'h10;
  assign mem[4989] = 5'h00;
  assign mem[4990] = 5'h01;
  assign mem[4991] = 5'h10;
  assign mem[4992] = 5'h00;
  assign mem[4993] = 5'h06;
  assign mem[4994] = 5'h15;
  assign mem[4995] = 5'h14;
  assign mem[4996] = 5'h13;
  assign mem[4997] = 5'h12;
  assign mem[4998] = 5'h11;
  assign mem[4999] = 5'h10;
  assign mem[5000] = 5'h00;
  assign mem[5001] = 5'h01;
  assign mem[5002] = 5'h10;
  assign mem[5003] = 5'h00;
  assign mem[5004] = 5'h02;
  assign mem[5005] = 5'h11;
  assign mem[5006] = 5'h10;
  assign mem[5007] = 5'h00;
  assign mem[5008] = 5'h01;
  assign mem[5009] = 5'h10;
  assign mem[5010] = 5'h00;
  assign mem[5011] = 5'h03;
  assign mem[5012] = 5'h12;
  assign mem[5013] = 5'h11;
  assign mem[5014] = 5'h10;
  assign mem[5015] = 5'h00;
  assign mem[5016] = 5'h01;
  assign mem[5017] = 5'h10;
  assign mem[5018] = 5'h00;
  assign mem[5019] = 5'h02;
  assign mem[5020] = 5'h11;
  assign mem[5021] = 5'h10;
  assign mem[5022] = 5'h00;
  assign mem[5023] = 5'h01;
  assign mem[5024] = 5'h10;
  assign mem[5025] = 5'h00;
  assign mem[5026] = 5'h04;
  assign mem[5027] = 5'h13;
  assign mem[5028] = 5'h12;
  assign mem[5029] = 5'h11;
  assign mem[5030] = 5'h10;
  assign mem[5031] = 5'h00;
  assign mem[5032] = 5'h01;
  assign mem[5033] = 5'h10;
  assign mem[5034] = 5'h00;
  assign mem[5035] = 5'h02;
  assign mem[5036] = 5'h11;
  assign mem[5037] = 5'h10;
  assign mem[5038] = 5'h00;
  assign mem[5039] = 5'h01;
  assign mem[5040] = 5'h10;
  assign mem[5041] = 5'h00;
  assign mem[5042] = 5'h03;
  assign mem[5043] = 5'h12;
  assign mem[5044] = 5'h11;
  assign mem[5045] = 5'h10;
  assign mem[5046] = 5'h00;
  assign mem[5047] = 5'h01;
  assign mem[5048] = 5'h10;
  assign mem[5049] = 5'h00;
  assign mem[5050] = 5'h02;
  assign mem[5051] = 5'h11;
  assign mem[5052] = 5'h10;
  assign mem[5053] = 5'h00;
  assign mem[5054] = 5'h01;
  assign mem[5055] = 5'h10;
  assign mem[5056] = 5'h00;
  assign mem[5057] = 5'h05;
  assign mem[5058] = 5'h14;
  assign mem[5059] = 5'h13;
  assign mem[5060] = 5'h12;
  assign mem[5061] = 5'h11;
  assign mem[5062] = 5'h10;
  assign mem[5063] = 5'h00;
  assign mem[5064] = 5'h01;
  assign mem[5065] = 5'h10;
  assign mem[5066] = 5'h00;
  assign mem[5067] = 5'h02;
  assign mem[5068] = 5'h11;
  assign mem[5069] = 5'h10;
  assign mem[5070] = 5'h00;
  assign mem[5071] = 5'h01;
  assign mem[5072] = 5'h10;
  assign mem[5073] = 5'h00;
  assign mem[5074] = 5'h03;
  assign mem[5075] = 5'h12;
  assign mem[5076] = 5'h11;
  assign mem[5077] = 5'h10;
  assign mem[5078] = 5'h00;
  assign mem[5079] = 5'h01;
  assign mem[5080] = 5'h10;
  assign mem[5081] = 5'h00;
  assign mem[5082] = 5'h02;
  assign mem[5083] = 5'h11;
  assign mem[5084] = 5'h10;
  assign mem[5085] = 5'h00;
  assign mem[5086] = 5'h01;
  assign mem[5087] = 5'h10;
  assign mem[5088] = 5'h00;
  assign mem[5089] = 5'h04;
  assign mem[5090] = 5'h13;
  assign mem[5091] = 5'h12;
  assign mem[5092] = 5'h11;
  assign mem[5093] = 5'h10;
  assign mem[5094] = 5'h00;
  assign mem[5095] = 5'h01;
  assign mem[5096] = 5'h10;
  assign mem[5097] = 5'h00;
  assign mem[5098] = 5'h02;
  assign mem[5099] = 5'h11;
  assign mem[5100] = 5'h10;
  assign mem[5101] = 5'h00;
  assign mem[5102] = 5'h01;
  assign mem[5103] = 5'h10;
  assign mem[5104] = 5'h00;
  assign mem[5105] = 5'h03;
  assign mem[5106] = 5'h12;
  assign mem[5107] = 5'h11;
  assign mem[5108] = 5'h10;
  assign mem[5109] = 5'h00;
  assign mem[5110] = 5'h01;
  assign mem[5111] = 5'h10;
  assign mem[5112] = 5'h00;
  assign mem[5113] = 5'h02;
  assign mem[5114] = 5'h11;
  assign mem[5115] = 5'h10;
  assign mem[5116] = 5'h00;
  assign mem[5117] = 5'h01;
  assign mem[5118] = 5'h10;
  assign mem[5119] = 5'h00;
  assign mem[5120] = 5'h09;
  assign mem[5121] = 5'h18;
  assign mem[5122] = 5'h17;
  assign mem[5123] = 5'h16;
  assign mem[5124] = 5'h15;
  assign mem[5125] = 5'h14;
  assign mem[5126] = 5'h13;
  assign mem[5127] = 5'h12;
  assign mem[5128] = 5'h11;
  assign mem[5129] = 5'h10;
  assign mem[5130] = 5'h00;
  assign mem[5131] = 5'h01;
  assign mem[5132] = 5'h10;
  assign mem[5133] = 5'h00;
  assign mem[5134] = 5'h02;
  assign mem[5135] = 5'h11;
  assign mem[5136] = 5'h10;
  assign mem[5137] = 5'h00;
  assign mem[5138] = 5'h01;
  assign mem[5139] = 5'h10;
  assign mem[5140] = 5'h00;
  assign mem[5141] = 5'h03;
  assign mem[5142] = 5'h12;
  assign mem[5143] = 5'h11;
  assign mem[5144] = 5'h10;
  assign mem[5145] = 5'h00;
  assign mem[5146] = 5'h01;
  assign mem[5147] = 5'h10;
  assign mem[5148] = 5'h00;
  assign mem[5149] = 5'h02;
  assign mem[5150] = 5'h11;
  assign mem[5151] = 5'h10;
  assign mem[5152] = 5'h00;
  assign mem[5153] = 5'h01;
  assign mem[5154] = 5'h10;
  assign mem[5155] = 5'h00;
  assign mem[5156] = 5'h04;
  assign mem[5157] = 5'h13;
  assign mem[5158] = 5'h12;
  assign mem[5159] = 5'h11;
  assign mem[5160] = 5'h10;
  assign mem[5161] = 5'h00;
  assign mem[5162] = 5'h01;
  assign mem[5163] = 5'h10;
  assign mem[5164] = 5'h00;
  assign mem[5165] = 5'h02;
  assign mem[5166] = 5'h11;
  assign mem[5167] = 5'h10;
  assign mem[5168] = 5'h00;
  assign mem[5169] = 5'h01;
  assign mem[5170] = 5'h10;
  assign mem[5171] = 5'h00;
  assign mem[5172] = 5'h03;
  assign mem[5173] = 5'h12;
  assign mem[5174] = 5'h11;
  assign mem[5175] = 5'h10;
  assign mem[5176] = 5'h00;
  assign mem[5177] = 5'h01;
  assign mem[5178] = 5'h10;
  assign mem[5179] = 5'h00;
  assign mem[5180] = 5'h02;
  assign mem[5181] = 5'h11;
  assign mem[5182] = 5'h10;
  assign mem[5183] = 5'h00;
  assign mem[5184] = 5'h01;
  assign mem[5185] = 5'h10;
  assign mem[5186] = 5'h00;
  assign mem[5187] = 5'h05;
  assign mem[5188] = 5'h14;
  assign mem[5189] = 5'h13;
  assign mem[5190] = 5'h12;
  assign mem[5191] = 5'h11;
  assign mem[5192] = 5'h10;
  assign mem[5193] = 5'h00;
  assign mem[5194] = 5'h01;
  assign mem[5195] = 5'h10;
  assign mem[5196] = 5'h00;
  assign mem[5197] = 5'h02;
  assign mem[5198] = 5'h11;
  assign mem[5199] = 5'h10;
  assign mem[5200] = 5'h00;
  assign mem[5201] = 5'h01;
  assign mem[5202] = 5'h10;
  assign mem[5203] = 5'h00;
  assign mem[5204] = 5'h03;
  assign mem[5205] = 5'h12;
  assign mem[5206] = 5'h11;
  assign mem[5207] = 5'h10;
  assign mem[5208] = 5'h00;
  assign mem[5209] = 5'h01;
  assign mem[5210] = 5'h10;
  assign mem[5211] = 5'h00;
  assign mem[5212] = 5'h02;
  assign mem[5213] = 5'h11;
  assign mem[5214] = 5'h10;
  assign mem[5215] = 5'h00;
  assign mem[5216] = 5'h01;
  assign mem[5217] = 5'h10;
  assign mem[5218] = 5'h00;
  assign mem[5219] = 5'h04;
  assign mem[5220] = 5'h13;
  assign mem[5221] = 5'h12;
  assign mem[5222] = 5'h11;
  assign mem[5223] = 5'h10;
  assign mem[5224] = 5'h00;
  assign mem[5225] = 5'h01;
  assign mem[5226] = 5'h10;
  assign mem[5227] = 5'h00;
  assign mem[5228] = 5'h02;
  assign mem[5229] = 5'h11;
  assign mem[5230] = 5'h10;
  assign mem[5231] = 5'h00;
  assign mem[5232] = 5'h01;
  assign mem[5233] = 5'h10;
  assign mem[5234] = 5'h00;
  assign mem[5235] = 5'h03;
  assign mem[5236] = 5'h12;
  assign mem[5237] = 5'h11;
  assign mem[5238] = 5'h10;
  assign mem[5239] = 5'h00;
  assign mem[5240] = 5'h01;
  assign mem[5241] = 5'h10;
  assign mem[5242] = 5'h00;
  assign mem[5243] = 5'h02;
  assign mem[5244] = 5'h11;
  assign mem[5245] = 5'h10;
  assign mem[5246] = 5'h00;
  assign mem[5247] = 5'h01;
  assign mem[5248] = 5'h10;
  assign mem[5249] = 5'h00;
  assign mem[5250] = 5'h06;
  assign mem[5251] = 5'h15;
  assign mem[5252] = 5'h14;
  assign mem[5253] = 5'h13;
  assign mem[5254] = 5'h12;
  assign mem[5255] = 5'h11;
  assign mem[5256] = 5'h10;
  assign mem[5257] = 5'h00;
  assign mem[5258] = 5'h01;
  assign mem[5259] = 5'h10;
  assign mem[5260] = 5'h00;
  assign mem[5261] = 5'h02;
  assign mem[5262] = 5'h11;
  assign mem[5263] = 5'h10;
  assign mem[5264] = 5'h00;
  assign mem[5265] = 5'h01;
  assign mem[5266] = 5'h10;
  assign mem[5267] = 5'h00;
  assign mem[5268] = 5'h03;
  assign mem[5269] = 5'h12;
  assign mem[5270] = 5'h11;
  assign mem[5271] = 5'h10;
  assign mem[5272] = 5'h00;
  assign mem[5273] = 5'h01;
  assign mem[5274] = 5'h10;
  assign mem[5275] = 5'h00;
  assign mem[5276] = 5'h02;
  assign mem[5277] = 5'h11;
  assign mem[5278] = 5'h10;
  assign mem[5279] = 5'h00;
  assign mem[5280] = 5'h01;
  assign mem[5281] = 5'h10;
  assign mem[5282] = 5'h00;
  assign mem[5283] = 5'h04;
  assign mem[5284] = 5'h13;
  assign mem[5285] = 5'h12;
  assign mem[5286] = 5'h11;
  assign mem[5287] = 5'h10;
  assign mem[5288] = 5'h00;
  assign mem[5289] = 5'h01;
  assign mem[5290] = 5'h10;
  assign mem[5291] = 5'h00;
  assign mem[5292] = 5'h02;
  assign mem[5293] = 5'h11;
  assign mem[5294] = 5'h10;
  assign mem[5295] = 5'h00;
  assign mem[5296] = 5'h01;
  assign mem[5297] = 5'h10;
  assign mem[5298] = 5'h00;
  assign mem[5299] = 5'h03;
  assign mem[5300] = 5'h12;
  assign mem[5301] = 5'h11;
  assign mem[5302] = 5'h10;
  assign mem[5303] = 5'h00;
  assign mem[5304] = 5'h01;
  assign mem[5305] = 5'h10;
  assign mem[5306] = 5'h00;
  assign mem[5307] = 5'h02;
  assign mem[5308] = 5'h11;
  assign mem[5309] = 5'h10;
  assign mem[5310] = 5'h00;
  assign mem[5311] = 5'h01;
  assign mem[5312] = 5'h10;
  assign mem[5313] = 5'h00;
  assign mem[5314] = 5'h05;
  assign mem[5315] = 5'h14;
  assign mem[5316] = 5'h13;
  assign mem[5317] = 5'h12;
  assign mem[5318] = 5'h11;
  assign mem[5319] = 5'h10;
  assign mem[5320] = 5'h00;
  assign mem[5321] = 5'h01;
  assign mem[5322] = 5'h10;
  assign mem[5323] = 5'h00;
  assign mem[5324] = 5'h02;
  assign mem[5325] = 5'h11;
  assign mem[5326] = 5'h10;
  assign mem[5327] = 5'h00;
  assign mem[5328] = 5'h01;
  assign mem[5329] = 5'h10;
  assign mem[5330] = 5'h00;
  assign mem[5331] = 5'h03;
  assign mem[5332] = 5'h12;
  assign mem[5333] = 5'h11;
  assign mem[5334] = 5'h10;
  assign mem[5335] = 5'h00;
  assign mem[5336] = 5'h01;
  assign mem[5337] = 5'h10;
  assign mem[5338] = 5'h00;
  assign mem[5339] = 5'h02;
  assign mem[5340] = 5'h11;
  assign mem[5341] = 5'h10;
  assign mem[5342] = 5'h00;
  assign mem[5343] = 5'h01;
  assign mem[5344] = 5'h10;
  assign mem[5345] = 5'h00;
  assign mem[5346] = 5'h04;
  assign mem[5347] = 5'h13;
  assign mem[5348] = 5'h12;
  assign mem[5349] = 5'h11;
  assign mem[5350] = 5'h10;
  assign mem[5351] = 5'h00;
  assign mem[5352] = 5'h01;
  assign mem[5353] = 5'h10;
  assign mem[5354] = 5'h00;
  assign mem[5355] = 5'h02;
  assign mem[5356] = 5'h11;
  assign mem[5357] = 5'h10;
  assign mem[5358] = 5'h00;
  assign mem[5359] = 5'h01;
  assign mem[5360] = 5'h10;
  assign mem[5361] = 5'h00;
  assign mem[5362] = 5'h03;
  assign mem[5363] = 5'h12;
  assign mem[5364] = 5'h11;
  assign mem[5365] = 5'h10;
  assign mem[5366] = 5'h00;
  assign mem[5367] = 5'h01;
  assign mem[5368] = 5'h10;
  assign mem[5369] = 5'h00;
  assign mem[5370] = 5'h02;
  assign mem[5371] = 5'h11;
  assign mem[5372] = 5'h10;
  assign mem[5373] = 5'h00;
  assign mem[5374] = 5'h01;
  assign mem[5375] = 5'h10;
  assign mem[5376] = 5'h00;
  assign mem[5377] = 5'h07;
  assign mem[5378] = 5'h16;
  assign mem[5379] = 5'h15;
  assign mem[5380] = 5'h14;
  assign mem[5381] = 5'h13;
  assign mem[5382] = 5'h12;
  assign mem[5383] = 5'h11;
  assign mem[5384] = 5'h10;
  assign mem[5385] = 5'h00;
  assign mem[5386] = 5'h01;
  assign mem[5387] = 5'h10;
  assign mem[5388] = 5'h00;
  assign mem[5389] = 5'h02;
  assign mem[5390] = 5'h11;
  assign mem[5391] = 5'h10;
  assign mem[5392] = 5'h00;
  assign mem[5393] = 5'h01;
  assign mem[5394] = 5'h10;
  assign mem[5395] = 5'h00;
  assign mem[5396] = 5'h03;
  assign mem[5397] = 5'h12;
  assign mem[5398] = 5'h11;
  assign mem[5399] = 5'h10;
  assign mem[5400] = 5'h00;
  assign mem[5401] = 5'h01;
  assign mem[5402] = 5'h10;
  assign mem[5403] = 5'h00;
  assign mem[5404] = 5'h02;
  assign mem[5405] = 5'h11;
  assign mem[5406] = 5'h10;
  assign mem[5407] = 5'h00;
  assign mem[5408] = 5'h01;
  assign mem[5409] = 5'h10;
  assign mem[5410] = 5'h00;
  assign mem[5411] = 5'h04;
  assign mem[5412] = 5'h13;
  assign mem[5413] = 5'h12;
  assign mem[5414] = 5'h11;
  assign mem[5415] = 5'h10;
  assign mem[5416] = 5'h00;
  assign mem[5417] = 5'h01;
  assign mem[5418] = 5'h10;
  assign mem[5419] = 5'h00;
  assign mem[5420] = 5'h02;
  assign mem[5421] = 5'h11;
  assign mem[5422] = 5'h10;
  assign mem[5423] = 5'h00;
  assign mem[5424] = 5'h01;
  assign mem[5425] = 5'h10;
  assign mem[5426] = 5'h00;
  assign mem[5427] = 5'h03;
  assign mem[5428] = 5'h12;
  assign mem[5429] = 5'h11;
  assign mem[5430] = 5'h10;
  assign mem[5431] = 5'h00;
  assign mem[5432] = 5'h01;
  assign mem[5433] = 5'h10;
  assign mem[5434] = 5'h00;
  assign mem[5435] = 5'h02;
  assign mem[5436] = 5'h11;
  assign mem[5437] = 5'h10;
  assign mem[5438] = 5'h00;
  assign mem[5439] = 5'h01;
  assign mem[5440] = 5'h10;
  assign mem[5441] = 5'h00;
  assign mem[5442] = 5'h05;
  assign mem[5443] = 5'h14;
  assign mem[5444] = 5'h13;
  assign mem[5445] = 5'h12;
  assign mem[5446] = 5'h11;
  assign mem[5447] = 5'h10;
  assign mem[5448] = 5'h00;
  assign mem[5449] = 5'h01;
  assign mem[5450] = 5'h10;
  assign mem[5451] = 5'h00;
  assign mem[5452] = 5'h02;
  assign mem[5453] = 5'h11;
  assign mem[5454] = 5'h10;
  assign mem[5455] = 5'h00;
  assign mem[5456] = 5'h01;
  assign mem[5457] = 5'h10;
  assign mem[5458] = 5'h00;
  assign mem[5459] = 5'h03;
  assign mem[5460] = 5'h12;
  assign mem[5461] = 5'h11;
  assign mem[5462] = 5'h10;
  assign mem[5463] = 5'h00;
  assign mem[5464] = 5'h01;
  assign mem[5465] = 5'h10;
  assign mem[5466] = 5'h00;
  assign mem[5467] = 5'h02;
  assign mem[5468] = 5'h11;
  assign mem[5469] = 5'h10;
  assign mem[5470] = 5'h00;
  assign mem[5471] = 5'h01;
  assign mem[5472] = 5'h10;
  assign mem[5473] = 5'h00;
  assign mem[5474] = 5'h04;
  assign mem[5475] = 5'h13;
  assign mem[5476] = 5'h12;
  assign mem[5477] = 5'h11;
  assign mem[5478] = 5'h10;
  assign mem[5479] = 5'h00;
  assign mem[5480] = 5'h01;
  assign mem[5481] = 5'h10;
  assign mem[5482] = 5'h00;
  assign mem[5483] = 5'h02;
  assign mem[5484] = 5'h11;
  assign mem[5485] = 5'h10;
  assign mem[5486] = 5'h00;
  assign mem[5487] = 5'h01;
  assign mem[5488] = 5'h10;
  assign mem[5489] = 5'h00;
  assign mem[5490] = 5'h03;
  assign mem[5491] = 5'h12;
  assign mem[5492] = 5'h11;
  assign mem[5493] = 5'h10;
  assign mem[5494] = 5'h00;
  assign mem[5495] = 5'h01;
  assign mem[5496] = 5'h10;
  assign mem[5497] = 5'h00;
  assign mem[5498] = 5'h02;
  assign mem[5499] = 5'h11;
  assign mem[5500] = 5'h10;
  assign mem[5501] = 5'h00;
  assign mem[5502] = 5'h01;
  assign mem[5503] = 5'h10;
  assign mem[5504] = 5'h00;
  assign mem[5505] = 5'h06;
  assign mem[5506] = 5'h15;
  assign mem[5507] = 5'h14;
  assign mem[5508] = 5'h13;
  assign mem[5509] = 5'h12;
  assign mem[5510] = 5'h11;
  assign mem[5511] = 5'h10;
  assign mem[5512] = 5'h00;
  assign mem[5513] = 5'h01;
  assign mem[5514] = 5'h10;
  assign mem[5515] = 5'h00;
  assign mem[5516] = 5'h02;
  assign mem[5517] = 5'h11;
  assign mem[5518] = 5'h10;
  assign mem[5519] = 5'h00;
  assign mem[5520] = 5'h01;
  assign mem[5521] = 5'h10;
  assign mem[5522] = 5'h00;
  assign mem[5523] = 5'h03;
  assign mem[5524] = 5'h12;
  assign mem[5525] = 5'h11;
  assign mem[5526] = 5'h10;
  assign mem[5527] = 5'h00;
  assign mem[5528] = 5'h01;
  assign mem[5529] = 5'h10;
  assign mem[5530] = 5'h00;
  assign mem[5531] = 5'h02;
  assign mem[5532] = 5'h11;
  assign mem[5533] = 5'h10;
  assign mem[5534] = 5'h00;
  assign mem[5535] = 5'h01;
  assign mem[5536] = 5'h10;
  assign mem[5537] = 5'h00;
  assign mem[5538] = 5'h04;
  assign mem[5539] = 5'h13;
  assign mem[5540] = 5'h12;
  assign mem[5541] = 5'h11;
  assign mem[5542] = 5'h10;
  assign mem[5543] = 5'h00;
  assign mem[5544] = 5'h01;
  assign mem[5545] = 5'h10;
  assign mem[5546] = 5'h00;
  assign mem[5547] = 5'h02;
  assign mem[5548] = 5'h11;
  assign mem[5549] = 5'h10;
  assign mem[5550] = 5'h00;
  assign mem[5551] = 5'h01;
  assign mem[5552] = 5'h10;
  assign mem[5553] = 5'h00;
  assign mem[5554] = 5'h03;
  assign mem[5555] = 5'h12;
  assign mem[5556] = 5'h11;
  assign mem[5557] = 5'h10;
  assign mem[5558] = 5'h00;
  assign mem[5559] = 5'h01;
  assign mem[5560] = 5'h10;
  assign mem[5561] = 5'h00;
  assign mem[5562] = 5'h02;
  assign mem[5563] = 5'h11;
  assign mem[5564] = 5'h10;
  assign mem[5565] = 5'h00;
  assign mem[5566] = 5'h01;
  assign mem[5567] = 5'h10;
  assign mem[5568] = 5'h00;
  assign mem[5569] = 5'h05;
  assign mem[5570] = 5'h14;
  assign mem[5571] = 5'h13;
  assign mem[5572] = 5'h12;
  assign mem[5573] = 5'h11;
  assign mem[5574] = 5'h10;
  assign mem[5575] = 5'h00;
  assign mem[5576] = 5'h01;
  assign mem[5577] = 5'h10;
  assign mem[5578] = 5'h00;
  assign mem[5579] = 5'h02;
  assign mem[5580] = 5'h11;
  assign mem[5581] = 5'h10;
  assign mem[5582] = 5'h00;
  assign mem[5583] = 5'h01;
  assign mem[5584] = 5'h10;
  assign mem[5585] = 5'h00;
  assign mem[5586] = 5'h03;
  assign mem[5587] = 5'h12;
  assign mem[5588] = 5'h11;
  assign mem[5589] = 5'h10;
  assign mem[5590] = 5'h00;
  assign mem[5591] = 5'h01;
  assign mem[5592] = 5'h10;
  assign mem[5593] = 5'h00;
  assign mem[5594] = 5'h02;
  assign mem[5595] = 5'h11;
  assign mem[5596] = 5'h10;
  assign mem[5597] = 5'h00;
  assign mem[5598] = 5'h01;
  assign mem[5599] = 5'h10;
  assign mem[5600] = 5'h00;
  assign mem[5601] = 5'h04;
  assign mem[5602] = 5'h13;
  assign mem[5603] = 5'h12;
  assign mem[5604] = 5'h11;
  assign mem[5605] = 5'h10;
  assign mem[5606] = 5'h00;
  assign mem[5607] = 5'h01;
  assign mem[5608] = 5'h10;
  assign mem[5609] = 5'h00;
  assign mem[5610] = 5'h02;
  assign mem[5611] = 5'h11;
  assign mem[5612] = 5'h10;
  assign mem[5613] = 5'h00;
  assign mem[5614] = 5'h01;
  assign mem[5615] = 5'h10;
  assign mem[5616] = 5'h00;
  assign mem[5617] = 5'h03;
  assign mem[5618] = 5'h12;
  assign mem[5619] = 5'h11;
  assign mem[5620] = 5'h10;
  assign mem[5621] = 5'h00;
  assign mem[5622] = 5'h01;
  assign mem[5623] = 5'h10;
  assign mem[5624] = 5'h00;
  assign mem[5625] = 5'h02;
  assign mem[5626] = 5'h11;
  assign mem[5627] = 5'h10;
  assign mem[5628] = 5'h00;
  assign mem[5629] = 5'h01;
  assign mem[5630] = 5'h10;
  assign mem[5631] = 5'h00;
  assign mem[5632] = 5'h08;
  assign mem[5633] = 5'h17;
  assign mem[5634] = 5'h16;
  assign mem[5635] = 5'h15;
  assign mem[5636] = 5'h14;
  assign mem[5637] = 5'h13;
  assign mem[5638] = 5'h12;
  assign mem[5639] = 5'h11;
  assign mem[5640] = 5'h10;
  assign mem[5641] = 5'h00;
  assign mem[5642] = 5'h01;
  assign mem[5643] = 5'h10;
  assign mem[5644] = 5'h00;
  assign mem[5645] = 5'h02;
  assign mem[5646] = 5'h11;
  assign mem[5647] = 5'h10;
  assign mem[5648] = 5'h00;
  assign mem[5649] = 5'h01;
  assign mem[5650] = 5'h10;
  assign mem[5651] = 5'h00;
  assign mem[5652] = 5'h03;
  assign mem[5653] = 5'h12;
  assign mem[5654] = 5'h11;
  assign mem[5655] = 5'h10;
  assign mem[5656] = 5'h00;
  assign mem[5657] = 5'h01;
  assign mem[5658] = 5'h10;
  assign mem[5659] = 5'h00;
  assign mem[5660] = 5'h02;
  assign mem[5661] = 5'h11;
  assign mem[5662] = 5'h10;
  assign mem[5663] = 5'h00;
  assign mem[5664] = 5'h01;
  assign mem[5665] = 5'h10;
  assign mem[5666] = 5'h00;
  assign mem[5667] = 5'h04;
  assign mem[5668] = 5'h13;
  assign mem[5669] = 5'h12;
  assign mem[5670] = 5'h11;
  assign mem[5671] = 5'h10;
  assign mem[5672] = 5'h00;
  assign mem[5673] = 5'h01;
  assign mem[5674] = 5'h10;
  assign mem[5675] = 5'h00;
  assign mem[5676] = 5'h02;
  assign mem[5677] = 5'h11;
  assign mem[5678] = 5'h10;
  assign mem[5679] = 5'h00;
  assign mem[5680] = 5'h01;
  assign mem[5681] = 5'h10;
  assign mem[5682] = 5'h00;
  assign mem[5683] = 5'h03;
  assign mem[5684] = 5'h12;
  assign mem[5685] = 5'h11;
  assign mem[5686] = 5'h10;
  assign mem[5687] = 5'h00;
  assign mem[5688] = 5'h01;
  assign mem[5689] = 5'h10;
  assign mem[5690] = 5'h00;
  assign mem[5691] = 5'h02;
  assign mem[5692] = 5'h11;
  assign mem[5693] = 5'h10;
  assign mem[5694] = 5'h00;
  assign mem[5695] = 5'h01;
  assign mem[5696] = 5'h10;
  assign mem[5697] = 5'h00;
  assign mem[5698] = 5'h05;
  assign mem[5699] = 5'h14;
  assign mem[5700] = 5'h13;
  assign mem[5701] = 5'h12;
  assign mem[5702] = 5'h11;
  assign mem[5703] = 5'h10;
  assign mem[5704] = 5'h00;
  assign mem[5705] = 5'h01;
  assign mem[5706] = 5'h10;
  assign mem[5707] = 5'h00;
  assign mem[5708] = 5'h02;
  assign mem[5709] = 5'h11;
  assign mem[5710] = 5'h10;
  assign mem[5711] = 5'h00;
  assign mem[5712] = 5'h01;
  assign mem[5713] = 5'h10;
  assign mem[5714] = 5'h00;
  assign mem[5715] = 5'h03;
  assign mem[5716] = 5'h12;
  assign mem[5717] = 5'h11;
  assign mem[5718] = 5'h10;
  assign mem[5719] = 5'h00;
  assign mem[5720] = 5'h01;
  assign mem[5721] = 5'h10;
  assign mem[5722] = 5'h00;
  assign mem[5723] = 5'h02;
  assign mem[5724] = 5'h11;
  assign mem[5725] = 5'h10;
  assign mem[5726] = 5'h00;
  assign mem[5727] = 5'h01;
  assign mem[5728] = 5'h10;
  assign mem[5729] = 5'h00;
  assign mem[5730] = 5'h04;
  assign mem[5731] = 5'h13;
  assign mem[5732] = 5'h12;
  assign mem[5733] = 5'h11;
  assign mem[5734] = 5'h10;
  assign mem[5735] = 5'h00;
  assign mem[5736] = 5'h01;
  assign mem[5737] = 5'h10;
  assign mem[5738] = 5'h00;
  assign mem[5739] = 5'h02;
  assign mem[5740] = 5'h11;
  assign mem[5741] = 5'h10;
  assign mem[5742] = 5'h00;
  assign mem[5743] = 5'h01;
  assign mem[5744] = 5'h10;
  assign mem[5745] = 5'h00;
  assign mem[5746] = 5'h03;
  assign mem[5747] = 5'h12;
  assign mem[5748] = 5'h11;
  assign mem[5749] = 5'h10;
  assign mem[5750] = 5'h00;
  assign mem[5751] = 5'h01;
  assign mem[5752] = 5'h10;
  assign mem[5753] = 5'h00;
  assign mem[5754] = 5'h02;
  assign mem[5755] = 5'h11;
  assign mem[5756] = 5'h10;
  assign mem[5757] = 5'h00;
  assign mem[5758] = 5'h01;
  assign mem[5759] = 5'h10;
  assign mem[5760] = 5'h00;
  assign mem[5761] = 5'h06;
  assign mem[5762] = 5'h15;
  assign mem[5763] = 5'h14;
  assign mem[5764] = 5'h13;
  assign mem[5765] = 5'h12;
  assign mem[5766] = 5'h11;
  assign mem[5767] = 5'h10;
  assign mem[5768] = 5'h00;
  assign mem[5769] = 5'h01;
  assign mem[5770] = 5'h10;
  assign mem[5771] = 5'h00;
  assign mem[5772] = 5'h02;
  assign mem[5773] = 5'h11;
  assign mem[5774] = 5'h10;
  assign mem[5775] = 5'h00;
  assign mem[5776] = 5'h01;
  assign mem[5777] = 5'h10;
  assign mem[5778] = 5'h00;
  assign mem[5779] = 5'h03;
  assign mem[5780] = 5'h12;
  assign mem[5781] = 5'h11;
  assign mem[5782] = 5'h10;
  assign mem[5783] = 5'h00;
  assign mem[5784] = 5'h01;
  assign mem[5785] = 5'h10;
  assign mem[5786] = 5'h00;
  assign mem[5787] = 5'h02;
  assign mem[5788] = 5'h11;
  assign mem[5789] = 5'h10;
  assign mem[5790] = 5'h00;
  assign mem[5791] = 5'h01;
  assign mem[5792] = 5'h10;
  assign mem[5793] = 5'h00;
  assign mem[5794] = 5'h04;
  assign mem[5795] = 5'h13;
  assign mem[5796] = 5'h12;
  assign mem[5797] = 5'h11;
  assign mem[5798] = 5'h10;
  assign mem[5799] = 5'h00;
  assign mem[5800] = 5'h01;
  assign mem[5801] = 5'h10;
  assign mem[5802] = 5'h00;
  assign mem[5803] = 5'h02;
  assign mem[5804] = 5'h11;
  assign mem[5805] = 5'h10;
  assign mem[5806] = 5'h00;
  assign mem[5807] = 5'h01;
  assign mem[5808] = 5'h10;
  assign mem[5809] = 5'h00;
  assign mem[5810] = 5'h03;
  assign mem[5811] = 5'h12;
  assign mem[5812] = 5'h11;
  assign mem[5813] = 5'h10;
  assign mem[5814] = 5'h00;
  assign mem[5815] = 5'h01;
  assign mem[5816] = 5'h10;
  assign mem[5817] = 5'h00;
  assign mem[5818] = 5'h02;
  assign mem[5819] = 5'h11;
  assign mem[5820] = 5'h10;
  assign mem[5821] = 5'h00;
  assign mem[5822] = 5'h01;
  assign mem[5823] = 5'h10;
  assign mem[5824] = 5'h00;
  assign mem[5825] = 5'h05;
  assign mem[5826] = 5'h14;
  assign mem[5827] = 5'h13;
  assign mem[5828] = 5'h12;
  assign mem[5829] = 5'h11;
  assign mem[5830] = 5'h10;
  assign mem[5831] = 5'h00;
  assign mem[5832] = 5'h01;
  assign mem[5833] = 5'h10;
  assign mem[5834] = 5'h00;
  assign mem[5835] = 5'h02;
  assign mem[5836] = 5'h11;
  assign mem[5837] = 5'h10;
  assign mem[5838] = 5'h00;
  assign mem[5839] = 5'h01;
  assign mem[5840] = 5'h10;
  assign mem[5841] = 5'h00;
  assign mem[5842] = 5'h03;
  assign mem[5843] = 5'h12;
  assign mem[5844] = 5'h11;
  assign mem[5845] = 5'h10;
  assign mem[5846] = 5'h00;
  assign mem[5847] = 5'h01;
  assign mem[5848] = 5'h10;
  assign mem[5849] = 5'h00;
  assign mem[5850] = 5'h02;
  assign mem[5851] = 5'h11;
  assign mem[5852] = 5'h10;
  assign mem[5853] = 5'h00;
  assign mem[5854] = 5'h01;
  assign mem[5855] = 5'h10;
  assign mem[5856] = 5'h00;
  assign mem[5857] = 5'h04;
  assign mem[5858] = 5'h13;
  assign mem[5859] = 5'h12;
  assign mem[5860] = 5'h11;
  assign mem[5861] = 5'h10;
  assign mem[5862] = 5'h00;
  assign mem[5863] = 5'h01;
  assign mem[5864] = 5'h10;
  assign mem[5865] = 5'h00;
  assign mem[5866] = 5'h02;
  assign mem[5867] = 5'h11;
  assign mem[5868] = 5'h10;
  assign mem[5869] = 5'h00;
  assign mem[5870] = 5'h01;
  assign mem[5871] = 5'h10;
  assign mem[5872] = 5'h00;
  assign mem[5873] = 5'h03;
  assign mem[5874] = 5'h12;
  assign mem[5875] = 5'h11;
  assign mem[5876] = 5'h10;
  assign mem[5877] = 5'h00;
  assign mem[5878] = 5'h01;
  assign mem[5879] = 5'h10;
  assign mem[5880] = 5'h00;
  assign mem[5881] = 5'h02;
  assign mem[5882] = 5'h11;
  assign mem[5883] = 5'h10;
  assign mem[5884] = 5'h00;
  assign mem[5885] = 5'h01;
  assign mem[5886] = 5'h10;
  assign mem[5887] = 5'h00;
  assign mem[5888] = 5'h07;
  assign mem[5889] = 5'h16;
  assign mem[5890] = 5'h15;
  assign mem[5891] = 5'h14;
  assign mem[5892] = 5'h13;
  assign mem[5893] = 5'h12;
  assign mem[5894] = 5'h11;
  assign mem[5895] = 5'h10;
  assign mem[5896] = 5'h00;
  assign mem[5897] = 5'h01;
  assign mem[5898] = 5'h10;
  assign mem[5899] = 5'h00;
  assign mem[5900] = 5'h02;
  assign mem[5901] = 5'h11;
  assign mem[5902] = 5'h10;
  assign mem[5903] = 5'h00;
  assign mem[5904] = 5'h01;
  assign mem[5905] = 5'h10;
  assign mem[5906] = 5'h00;
  assign mem[5907] = 5'h03;
  assign mem[5908] = 5'h12;
  assign mem[5909] = 5'h11;
  assign mem[5910] = 5'h10;
  assign mem[5911] = 5'h00;
  assign mem[5912] = 5'h01;
  assign mem[5913] = 5'h10;
  assign mem[5914] = 5'h00;
  assign mem[5915] = 5'h02;
  assign mem[5916] = 5'h11;
  assign mem[5917] = 5'h10;
  assign mem[5918] = 5'h00;
  assign mem[5919] = 5'h01;
  assign mem[5920] = 5'h10;
  assign mem[5921] = 5'h00;
  assign mem[5922] = 5'h04;
  assign mem[5923] = 5'h13;
  assign mem[5924] = 5'h12;
  assign mem[5925] = 5'h11;
  assign mem[5926] = 5'h10;
  assign mem[5927] = 5'h00;
  assign mem[5928] = 5'h01;
  assign mem[5929] = 5'h10;
  assign mem[5930] = 5'h00;
  assign mem[5931] = 5'h02;
  assign mem[5932] = 5'h11;
  assign mem[5933] = 5'h10;
  assign mem[5934] = 5'h00;
  assign mem[5935] = 5'h01;
  assign mem[5936] = 5'h10;
  assign mem[5937] = 5'h00;
  assign mem[5938] = 5'h03;
  assign mem[5939] = 5'h12;
  assign mem[5940] = 5'h11;
  assign mem[5941] = 5'h10;
  assign mem[5942] = 5'h00;
  assign mem[5943] = 5'h01;
  assign mem[5944] = 5'h10;
  assign mem[5945] = 5'h00;
  assign mem[5946] = 5'h02;
  assign mem[5947] = 5'h11;
  assign mem[5948] = 5'h10;
  assign mem[5949] = 5'h00;
  assign mem[5950] = 5'h01;
  assign mem[5951] = 5'h10;
  assign mem[5952] = 5'h00;
  assign mem[5953] = 5'h05;
  assign mem[5954] = 5'h14;
  assign mem[5955] = 5'h13;
  assign mem[5956] = 5'h12;
  assign mem[5957] = 5'h11;
  assign mem[5958] = 5'h10;
  assign mem[5959] = 5'h00;
  assign mem[5960] = 5'h01;
  assign mem[5961] = 5'h10;
  assign mem[5962] = 5'h00;
  assign mem[5963] = 5'h02;
  assign mem[5964] = 5'h11;
  assign mem[5965] = 5'h10;
  assign mem[5966] = 5'h00;
  assign mem[5967] = 5'h01;
  assign mem[5968] = 5'h10;
  assign mem[5969] = 5'h00;
  assign mem[5970] = 5'h03;
  assign mem[5971] = 5'h12;
  assign mem[5972] = 5'h11;
  assign mem[5973] = 5'h10;
  assign mem[5974] = 5'h00;
  assign mem[5975] = 5'h01;
  assign mem[5976] = 5'h10;
  assign mem[5977] = 5'h00;
  assign mem[5978] = 5'h02;
  assign mem[5979] = 5'h11;
  assign mem[5980] = 5'h10;
  assign mem[5981] = 5'h00;
  assign mem[5982] = 5'h01;
  assign mem[5983] = 5'h10;
  assign mem[5984] = 5'h00;
  assign mem[5985] = 5'h04;
  assign mem[5986] = 5'h13;
  assign mem[5987] = 5'h12;
  assign mem[5988] = 5'h11;
  assign mem[5989] = 5'h10;
  assign mem[5990] = 5'h00;
  assign mem[5991] = 5'h01;
  assign mem[5992] = 5'h10;
  assign mem[5993] = 5'h00;
  assign mem[5994] = 5'h02;
  assign mem[5995] = 5'h11;
  assign mem[5996] = 5'h10;
  assign mem[5997] = 5'h00;
  assign mem[5998] = 5'h01;
  assign mem[5999] = 5'h10;
  assign mem[6000] = 5'h00;
  assign mem[6001] = 5'h03;
  assign mem[6002] = 5'h12;
  assign mem[6003] = 5'h11;
  assign mem[6004] = 5'h10;
  assign mem[6005] = 5'h00;
  assign mem[6006] = 5'h01;
  assign mem[6007] = 5'h10;
  assign mem[6008] = 5'h00;
  assign mem[6009] = 5'h02;
  assign mem[6010] = 5'h11;
  assign mem[6011] = 5'h10;
  assign mem[6012] = 5'h00;
  assign mem[6013] = 5'h01;
  assign mem[6014] = 5'h10;
  assign mem[6015] = 5'h00;
  assign mem[6016] = 5'h06;
  assign mem[6017] = 5'h15;
  assign mem[6018] = 5'h14;
  assign mem[6019] = 5'h13;
  assign mem[6020] = 5'h12;
  assign mem[6021] = 5'h11;
  assign mem[6022] = 5'h10;
  assign mem[6023] = 5'h00;
  assign mem[6024] = 5'h01;
  assign mem[6025] = 5'h10;
  assign mem[6026] = 5'h00;
  assign mem[6027] = 5'h02;
  assign mem[6028] = 5'h11;
  assign mem[6029] = 5'h10;
  assign mem[6030] = 5'h00;
  assign mem[6031] = 5'h01;
  assign mem[6032] = 5'h10;
  assign mem[6033] = 5'h00;
  assign mem[6034] = 5'h03;
  assign mem[6035] = 5'h12;
  assign mem[6036] = 5'h11;
  assign mem[6037] = 5'h10;
  assign mem[6038] = 5'h00;
  assign mem[6039] = 5'h01;
  assign mem[6040] = 5'h10;
  assign mem[6041] = 5'h00;
  assign mem[6042] = 5'h02;
  assign mem[6043] = 5'h11;
  assign mem[6044] = 5'h10;
  assign mem[6045] = 5'h00;
  assign mem[6046] = 5'h01;
  assign mem[6047] = 5'h10;
  assign mem[6048] = 5'h00;
  assign mem[6049] = 5'h04;
  assign mem[6050] = 5'h13;
  assign mem[6051] = 5'h12;
  assign mem[6052] = 5'h11;
  assign mem[6053] = 5'h10;
  assign mem[6054] = 5'h00;
  assign mem[6055] = 5'h01;
  assign mem[6056] = 5'h10;
  assign mem[6057] = 5'h00;
  assign mem[6058] = 5'h02;
  assign mem[6059] = 5'h11;
  assign mem[6060] = 5'h10;
  assign mem[6061] = 5'h00;
  assign mem[6062] = 5'h01;
  assign mem[6063] = 5'h10;
  assign mem[6064] = 5'h00;
  assign mem[6065] = 5'h03;
  assign mem[6066] = 5'h12;
  assign mem[6067] = 5'h11;
  assign mem[6068] = 5'h10;
  assign mem[6069] = 5'h00;
  assign mem[6070] = 5'h01;
  assign mem[6071] = 5'h10;
  assign mem[6072] = 5'h00;
  assign mem[6073] = 5'h02;
  assign mem[6074] = 5'h11;
  assign mem[6075] = 5'h10;
  assign mem[6076] = 5'h00;
  assign mem[6077] = 5'h01;
  assign mem[6078] = 5'h10;
  assign mem[6079] = 5'h00;
  assign mem[6080] = 5'h05;
  assign mem[6081] = 5'h14;
  assign mem[6082] = 5'h13;
  assign mem[6083] = 5'h12;
  assign mem[6084] = 5'h11;
  assign mem[6085] = 5'h10;
  assign mem[6086] = 5'h00;
  assign mem[6087] = 5'h01;
  assign mem[6088] = 5'h10;
  assign mem[6089] = 5'h00;
  assign mem[6090] = 5'h02;
  assign mem[6091] = 5'h11;
  assign mem[6092] = 5'h10;
  assign mem[6093] = 5'h00;
  assign mem[6094] = 5'h01;
  assign mem[6095] = 5'h10;
  assign mem[6096] = 5'h00;
  assign mem[6097] = 5'h03;
  assign mem[6098] = 5'h12;
  assign mem[6099] = 5'h11;
  assign mem[6100] = 5'h10;
  assign mem[6101] = 5'h00;
  assign mem[6102] = 5'h01;
  assign mem[6103] = 5'h10;
  assign mem[6104] = 5'h00;
  assign mem[6105] = 5'h02;
  assign mem[6106] = 5'h11;
  assign mem[6107] = 5'h10;
  assign mem[6108] = 5'h00;
  assign mem[6109] = 5'h01;
  assign mem[6110] = 5'h10;
  assign mem[6111] = 5'h00;
  assign mem[6112] = 5'h04;
  assign mem[6113] = 5'h13;
  assign mem[6114] = 5'h12;
  assign mem[6115] = 5'h11;
  assign mem[6116] = 5'h10;
  assign mem[6117] = 5'h00;
  assign mem[6118] = 5'h01;
  assign mem[6119] = 5'h10;
  assign mem[6120] = 5'h00;
  assign mem[6121] = 5'h02;
  assign mem[6122] = 5'h11;
  assign mem[6123] = 5'h10;
  assign mem[6124] = 5'h00;
  assign mem[6125] = 5'h01;
  assign mem[6126] = 5'h10;
  assign mem[6127] = 5'h00;
  assign mem[6128] = 5'h03;
  assign mem[6129] = 5'h12;
  assign mem[6130] = 5'h11;
  assign mem[6131] = 5'h10;
  assign mem[6132] = 5'h00;
  assign mem[6133] = 5'h01;
  assign mem[6134] = 5'h10;
  assign mem[6135] = 5'h00;
  assign mem[6136] = 5'h02;
  assign mem[6137] = 5'h11;
  assign mem[6138] = 5'h10;
  assign mem[6139] = 5'h00;
  assign mem[6140] = 5'h01;
  assign mem[6141] = 5'h10;
  assign mem[6142] = 5'h00;
  assign mem[6143] = 5'h0a;
  assign mem[6144] = 5'h19;
  assign mem[6145] = 5'h18;
  assign mem[6146] = 5'h17;
  assign mem[6147] = 5'h16;
  assign mem[6148] = 5'h15;
  assign mem[6149] = 5'h14;
  assign mem[6150] = 5'h13;
  assign mem[6151] = 5'h12;
  assign mem[6152] = 5'h11;
  assign mem[6153] = 5'h10;
  assign mem[6154] = 5'h00;
  assign mem[6155] = 5'h01;
  assign mem[6156] = 5'h10;
  assign mem[6157] = 5'h00;
  assign mem[6158] = 5'h02;
  assign mem[6159] = 5'h11;
  assign mem[6160] = 5'h10;
  assign mem[6161] = 5'h00;
  assign mem[6162] = 5'h01;
  assign mem[6163] = 5'h10;
  assign mem[6164] = 5'h00;
  assign mem[6165] = 5'h03;
  assign mem[6166] = 5'h12;
  assign mem[6167] = 5'h11;
  assign mem[6168] = 5'h10;
  assign mem[6169] = 5'h00;
  assign mem[6170] = 5'h01;
  assign mem[6171] = 5'h10;
  assign mem[6172] = 5'h00;
  assign mem[6173] = 5'h02;
  assign mem[6174] = 5'h11;
  assign mem[6175] = 5'h10;
  assign mem[6176] = 5'h00;
  assign mem[6177] = 5'h01;
  assign mem[6178] = 5'h10;
  assign mem[6179] = 5'h00;
  assign mem[6180] = 5'h04;
  assign mem[6181] = 5'h13;
  assign mem[6182] = 5'h12;
  assign mem[6183] = 5'h11;
  assign mem[6184] = 5'h10;
  assign mem[6185] = 5'h00;
  assign mem[6186] = 5'h01;
  assign mem[6187] = 5'h10;
  assign mem[6188] = 5'h00;
  assign mem[6189] = 5'h02;
  assign mem[6190] = 5'h11;
  assign mem[6191] = 5'h10;
  assign mem[6192] = 5'h00;
  assign mem[6193] = 5'h01;
  assign mem[6194] = 5'h10;
  assign mem[6195] = 5'h00;
  assign mem[6196] = 5'h03;
  assign mem[6197] = 5'h12;
  assign mem[6198] = 5'h11;
  assign mem[6199] = 5'h10;
  assign mem[6200] = 5'h00;
  assign mem[6201] = 5'h01;
  assign mem[6202] = 5'h10;
  assign mem[6203] = 5'h00;
  assign mem[6204] = 5'h02;
  assign mem[6205] = 5'h11;
  assign mem[6206] = 5'h10;
  assign mem[6207] = 5'h00;
  assign mem[6208] = 5'h01;
  assign mem[6209] = 5'h10;
  assign mem[6210] = 5'h00;
  assign mem[6211] = 5'h05;
  assign mem[6212] = 5'h14;
  assign mem[6213] = 5'h13;
  assign mem[6214] = 5'h12;
  assign mem[6215] = 5'h11;
  assign mem[6216] = 5'h10;
  assign mem[6217] = 5'h00;
  assign mem[6218] = 5'h01;
  assign mem[6219] = 5'h10;
  assign mem[6220] = 5'h00;
  assign mem[6221] = 5'h02;
  assign mem[6222] = 5'h11;
  assign mem[6223] = 5'h10;
  assign mem[6224] = 5'h00;
  assign mem[6225] = 5'h01;
  assign mem[6226] = 5'h10;
  assign mem[6227] = 5'h00;
  assign mem[6228] = 5'h03;
  assign mem[6229] = 5'h12;
  assign mem[6230] = 5'h11;
  assign mem[6231] = 5'h10;
  assign mem[6232] = 5'h00;
  assign mem[6233] = 5'h01;
  assign mem[6234] = 5'h10;
  assign mem[6235] = 5'h00;
  assign mem[6236] = 5'h02;
  assign mem[6237] = 5'h11;
  assign mem[6238] = 5'h10;
  assign mem[6239] = 5'h00;
  assign mem[6240] = 5'h01;
  assign mem[6241] = 5'h10;
  assign mem[6242] = 5'h00;
  assign mem[6243] = 5'h04;
  assign mem[6244] = 5'h13;
  assign mem[6245] = 5'h12;
  assign mem[6246] = 5'h11;
  assign mem[6247] = 5'h10;
  assign mem[6248] = 5'h00;
  assign mem[6249] = 5'h01;
  assign mem[6250] = 5'h10;
  assign mem[6251] = 5'h00;
  assign mem[6252] = 5'h02;
  assign mem[6253] = 5'h11;
  assign mem[6254] = 5'h10;
  assign mem[6255] = 5'h00;
  assign mem[6256] = 5'h01;
  assign mem[6257] = 5'h10;
  assign mem[6258] = 5'h00;
  assign mem[6259] = 5'h03;
  assign mem[6260] = 5'h12;
  assign mem[6261] = 5'h11;
  assign mem[6262] = 5'h10;
  assign mem[6263] = 5'h00;
  assign mem[6264] = 5'h01;
  assign mem[6265] = 5'h10;
  assign mem[6266] = 5'h00;
  assign mem[6267] = 5'h02;
  assign mem[6268] = 5'h11;
  assign mem[6269] = 5'h10;
  assign mem[6270] = 5'h00;
  assign mem[6271] = 5'h01;
  assign mem[6272] = 5'h10;
  assign mem[6273] = 5'h00;
  assign mem[6274] = 5'h06;
  assign mem[6275] = 5'h15;
  assign mem[6276] = 5'h14;
  assign mem[6277] = 5'h13;
  assign mem[6278] = 5'h12;
  assign mem[6279] = 5'h11;
  assign mem[6280] = 5'h10;
  assign mem[6281] = 5'h00;
  assign mem[6282] = 5'h01;
  assign mem[6283] = 5'h10;
  assign mem[6284] = 5'h00;
  assign mem[6285] = 5'h02;
  assign mem[6286] = 5'h11;
  assign mem[6287] = 5'h10;
  assign mem[6288] = 5'h00;
  assign mem[6289] = 5'h01;
  assign mem[6290] = 5'h10;
  assign mem[6291] = 5'h00;
  assign mem[6292] = 5'h03;
  assign mem[6293] = 5'h12;
  assign mem[6294] = 5'h11;
  assign mem[6295] = 5'h10;
  assign mem[6296] = 5'h00;
  assign mem[6297] = 5'h01;
  assign mem[6298] = 5'h10;
  assign mem[6299] = 5'h00;
  assign mem[6300] = 5'h02;
  assign mem[6301] = 5'h11;
  assign mem[6302] = 5'h10;
  assign mem[6303] = 5'h00;
  assign mem[6304] = 5'h01;
  assign mem[6305] = 5'h10;
  assign mem[6306] = 5'h00;
  assign mem[6307] = 5'h04;
  assign mem[6308] = 5'h13;
  assign mem[6309] = 5'h12;
  assign mem[6310] = 5'h11;
  assign mem[6311] = 5'h10;
  assign mem[6312] = 5'h00;
  assign mem[6313] = 5'h01;
  assign mem[6314] = 5'h10;
  assign mem[6315] = 5'h00;
  assign mem[6316] = 5'h02;
  assign mem[6317] = 5'h11;
  assign mem[6318] = 5'h10;
  assign mem[6319] = 5'h00;
  assign mem[6320] = 5'h01;
  assign mem[6321] = 5'h10;
  assign mem[6322] = 5'h00;
  assign mem[6323] = 5'h03;
  assign mem[6324] = 5'h12;
  assign mem[6325] = 5'h11;
  assign mem[6326] = 5'h10;
  assign mem[6327] = 5'h00;
  assign mem[6328] = 5'h01;
  assign mem[6329] = 5'h10;
  assign mem[6330] = 5'h00;
  assign mem[6331] = 5'h02;
  assign mem[6332] = 5'h11;
  assign mem[6333] = 5'h10;
  assign mem[6334] = 5'h00;
  assign mem[6335] = 5'h01;
  assign mem[6336] = 5'h10;
  assign mem[6337] = 5'h00;
  assign mem[6338] = 5'h05;
  assign mem[6339] = 5'h14;
  assign mem[6340] = 5'h13;
  assign mem[6341] = 5'h12;
  assign mem[6342] = 5'h11;
  assign mem[6343] = 5'h10;
  assign mem[6344] = 5'h00;
  assign mem[6345] = 5'h01;
  assign mem[6346] = 5'h10;
  assign mem[6347] = 5'h00;
  assign mem[6348] = 5'h02;
  assign mem[6349] = 5'h11;
  assign mem[6350] = 5'h10;
  assign mem[6351] = 5'h00;
  assign mem[6352] = 5'h01;
  assign mem[6353] = 5'h10;
  assign mem[6354] = 5'h00;
  assign mem[6355] = 5'h03;
  assign mem[6356] = 5'h12;
  assign mem[6357] = 5'h11;
  assign mem[6358] = 5'h10;
  assign mem[6359] = 5'h00;
  assign mem[6360] = 5'h01;
  assign mem[6361] = 5'h10;
  assign mem[6362] = 5'h00;
  assign mem[6363] = 5'h02;
  assign mem[6364] = 5'h11;
  assign mem[6365] = 5'h10;
  assign mem[6366] = 5'h00;
  assign mem[6367] = 5'h01;
  assign mem[6368] = 5'h10;
  assign mem[6369] = 5'h00;
  assign mem[6370] = 5'h04;
  assign mem[6371] = 5'h13;
  assign mem[6372] = 5'h12;
  assign mem[6373] = 5'h11;
  assign mem[6374] = 5'h10;
  assign mem[6375] = 5'h00;
  assign mem[6376] = 5'h01;
  assign mem[6377] = 5'h10;
  assign mem[6378] = 5'h00;
  assign mem[6379] = 5'h02;
  assign mem[6380] = 5'h11;
  assign mem[6381] = 5'h10;
  assign mem[6382] = 5'h00;
  assign mem[6383] = 5'h01;
  assign mem[6384] = 5'h10;
  assign mem[6385] = 5'h00;
  assign mem[6386] = 5'h03;
  assign mem[6387] = 5'h12;
  assign mem[6388] = 5'h11;
  assign mem[6389] = 5'h10;
  assign mem[6390] = 5'h00;
  assign mem[6391] = 5'h01;
  assign mem[6392] = 5'h10;
  assign mem[6393] = 5'h00;
  assign mem[6394] = 5'h02;
  assign mem[6395] = 5'h11;
  assign mem[6396] = 5'h10;
  assign mem[6397] = 5'h00;
  assign mem[6398] = 5'h01;
  assign mem[6399] = 5'h10;
  assign mem[6400] = 5'h00;
  assign mem[6401] = 5'h07;
  assign mem[6402] = 5'h16;
  assign mem[6403] = 5'h15;
  assign mem[6404] = 5'h14;
  assign mem[6405] = 5'h13;
  assign mem[6406] = 5'h12;
  assign mem[6407] = 5'h11;
  assign mem[6408] = 5'h10;
  assign mem[6409] = 5'h00;
  assign mem[6410] = 5'h01;
  assign mem[6411] = 5'h10;
  assign mem[6412] = 5'h00;
  assign mem[6413] = 5'h02;
  assign mem[6414] = 5'h11;
  assign mem[6415] = 5'h10;
  assign mem[6416] = 5'h00;
  assign mem[6417] = 5'h01;
  assign mem[6418] = 5'h10;
  assign mem[6419] = 5'h00;
  assign mem[6420] = 5'h03;
  assign mem[6421] = 5'h12;
  assign mem[6422] = 5'h11;
  assign mem[6423] = 5'h10;
  assign mem[6424] = 5'h00;
  assign mem[6425] = 5'h01;
  assign mem[6426] = 5'h10;
  assign mem[6427] = 5'h00;
  assign mem[6428] = 5'h02;
  assign mem[6429] = 5'h11;
  assign mem[6430] = 5'h10;
  assign mem[6431] = 5'h00;
  assign mem[6432] = 5'h01;
  assign mem[6433] = 5'h10;
  assign mem[6434] = 5'h00;
  assign mem[6435] = 5'h04;
  assign mem[6436] = 5'h13;
  assign mem[6437] = 5'h12;
  assign mem[6438] = 5'h11;
  assign mem[6439] = 5'h10;
  assign mem[6440] = 5'h00;
  assign mem[6441] = 5'h01;
  assign mem[6442] = 5'h10;
  assign mem[6443] = 5'h00;
  assign mem[6444] = 5'h02;
  assign mem[6445] = 5'h11;
  assign mem[6446] = 5'h10;
  assign mem[6447] = 5'h00;
  assign mem[6448] = 5'h01;
  assign mem[6449] = 5'h10;
  assign mem[6450] = 5'h00;
  assign mem[6451] = 5'h03;
  assign mem[6452] = 5'h12;
  assign mem[6453] = 5'h11;
  assign mem[6454] = 5'h10;
  assign mem[6455] = 5'h00;
  assign mem[6456] = 5'h01;
  assign mem[6457] = 5'h10;
  assign mem[6458] = 5'h00;
  assign mem[6459] = 5'h02;
  assign mem[6460] = 5'h11;
  assign mem[6461] = 5'h10;
  assign mem[6462] = 5'h00;
  assign mem[6463] = 5'h01;
  assign mem[6464] = 5'h10;
  assign mem[6465] = 5'h00;
  assign mem[6466] = 5'h05;
  assign mem[6467] = 5'h14;
  assign mem[6468] = 5'h13;
  assign mem[6469] = 5'h12;
  assign mem[6470] = 5'h11;
  assign mem[6471] = 5'h10;
  assign mem[6472] = 5'h00;
  assign mem[6473] = 5'h01;
  assign mem[6474] = 5'h10;
  assign mem[6475] = 5'h00;
  assign mem[6476] = 5'h02;
  assign mem[6477] = 5'h11;
  assign mem[6478] = 5'h10;
  assign mem[6479] = 5'h00;
  assign mem[6480] = 5'h01;
  assign mem[6481] = 5'h10;
  assign mem[6482] = 5'h00;
  assign mem[6483] = 5'h03;
  assign mem[6484] = 5'h12;
  assign mem[6485] = 5'h11;
  assign mem[6486] = 5'h10;
  assign mem[6487] = 5'h00;
  assign mem[6488] = 5'h01;
  assign mem[6489] = 5'h10;
  assign mem[6490] = 5'h00;
  assign mem[6491] = 5'h02;
  assign mem[6492] = 5'h11;
  assign mem[6493] = 5'h10;
  assign mem[6494] = 5'h00;
  assign mem[6495] = 5'h01;
  assign mem[6496] = 5'h10;
  assign mem[6497] = 5'h00;
  assign mem[6498] = 5'h04;
  assign mem[6499] = 5'h13;
  assign mem[6500] = 5'h12;
  assign mem[6501] = 5'h11;
  assign mem[6502] = 5'h10;
  assign mem[6503] = 5'h00;
  assign mem[6504] = 5'h01;
  assign mem[6505] = 5'h10;
  assign mem[6506] = 5'h00;
  assign mem[6507] = 5'h02;
  assign mem[6508] = 5'h11;
  assign mem[6509] = 5'h10;
  assign mem[6510] = 5'h00;
  assign mem[6511] = 5'h01;
  assign mem[6512] = 5'h10;
  assign mem[6513] = 5'h00;
  assign mem[6514] = 5'h03;
  assign mem[6515] = 5'h12;
  assign mem[6516] = 5'h11;
  assign mem[6517] = 5'h10;
  assign mem[6518] = 5'h00;
  assign mem[6519] = 5'h01;
  assign mem[6520] = 5'h10;
  assign mem[6521] = 5'h00;
  assign mem[6522] = 5'h02;
  assign mem[6523] = 5'h11;
  assign mem[6524] = 5'h10;
  assign mem[6525] = 5'h00;
  assign mem[6526] = 5'h01;
  assign mem[6527] = 5'h10;
  assign mem[6528] = 5'h00;
  assign mem[6529] = 5'h06;
  assign mem[6530] = 5'h15;
  assign mem[6531] = 5'h14;
  assign mem[6532] = 5'h13;
  assign mem[6533] = 5'h12;
  assign mem[6534] = 5'h11;
  assign mem[6535] = 5'h10;
  assign mem[6536] = 5'h00;
  assign mem[6537] = 5'h01;
  assign mem[6538] = 5'h10;
  assign mem[6539] = 5'h00;
  assign mem[6540] = 5'h02;
  assign mem[6541] = 5'h11;
  assign mem[6542] = 5'h10;
  assign mem[6543] = 5'h00;
  assign mem[6544] = 5'h01;
  assign mem[6545] = 5'h10;
  assign mem[6546] = 5'h00;
  assign mem[6547] = 5'h03;
  assign mem[6548] = 5'h12;
  assign mem[6549] = 5'h11;
  assign mem[6550] = 5'h10;
  assign mem[6551] = 5'h00;
  assign mem[6552] = 5'h01;
  assign mem[6553] = 5'h10;
  assign mem[6554] = 5'h00;
  assign mem[6555] = 5'h02;
  assign mem[6556] = 5'h11;
  assign mem[6557] = 5'h10;
  assign mem[6558] = 5'h00;
  assign mem[6559] = 5'h01;
  assign mem[6560] = 5'h10;
  assign mem[6561] = 5'h00;
  assign mem[6562] = 5'h04;
  assign mem[6563] = 5'h13;
  assign mem[6564] = 5'h12;
  assign mem[6565] = 5'h11;
  assign mem[6566] = 5'h10;
  assign mem[6567] = 5'h00;
  assign mem[6568] = 5'h01;
  assign mem[6569] = 5'h10;
  assign mem[6570] = 5'h00;
  assign mem[6571] = 5'h02;
  assign mem[6572] = 5'h11;
  assign mem[6573] = 5'h10;
  assign mem[6574] = 5'h00;
  assign mem[6575] = 5'h01;
  assign mem[6576] = 5'h10;
  assign mem[6577] = 5'h00;
  assign mem[6578] = 5'h03;
  assign mem[6579] = 5'h12;
  assign mem[6580] = 5'h11;
  assign mem[6581] = 5'h10;
  assign mem[6582] = 5'h00;
  assign mem[6583] = 5'h01;
  assign mem[6584] = 5'h10;
  assign mem[6585] = 5'h00;
  assign mem[6586] = 5'h02;
  assign mem[6587] = 5'h11;
  assign mem[6588] = 5'h10;
  assign mem[6589] = 5'h00;
  assign mem[6590] = 5'h01;
  assign mem[6591] = 5'h10;
  assign mem[6592] = 5'h00;
  assign mem[6593] = 5'h05;
  assign mem[6594] = 5'h14;
  assign mem[6595] = 5'h13;
  assign mem[6596] = 5'h12;
  assign mem[6597] = 5'h11;
  assign mem[6598] = 5'h10;
  assign mem[6599] = 5'h00;
  assign mem[6600] = 5'h01;
  assign mem[6601] = 5'h10;
  assign mem[6602] = 5'h00;
  assign mem[6603] = 5'h02;
  assign mem[6604] = 5'h11;
  assign mem[6605] = 5'h10;
  assign mem[6606] = 5'h00;
  assign mem[6607] = 5'h01;
  assign mem[6608] = 5'h10;
  assign mem[6609] = 5'h00;
  assign mem[6610] = 5'h03;
  assign mem[6611] = 5'h12;
  assign mem[6612] = 5'h11;
  assign mem[6613] = 5'h10;
  assign mem[6614] = 5'h00;
  assign mem[6615] = 5'h01;
  assign mem[6616] = 5'h10;
  assign mem[6617] = 5'h00;
  assign mem[6618] = 5'h02;
  assign mem[6619] = 5'h11;
  assign mem[6620] = 5'h10;
  assign mem[6621] = 5'h00;
  assign mem[6622] = 5'h01;
  assign mem[6623] = 5'h10;
  assign mem[6624] = 5'h00;
  assign mem[6625] = 5'h04;
  assign mem[6626] = 5'h13;
  assign mem[6627] = 5'h12;
  assign mem[6628] = 5'h11;
  assign mem[6629] = 5'h10;
  assign mem[6630] = 5'h00;
  assign mem[6631] = 5'h01;
  assign mem[6632] = 5'h10;
  assign mem[6633] = 5'h00;
  assign mem[6634] = 5'h02;
  assign mem[6635] = 5'h11;
  assign mem[6636] = 5'h10;
  assign mem[6637] = 5'h00;
  assign mem[6638] = 5'h01;
  assign mem[6639] = 5'h10;
  assign mem[6640] = 5'h00;
  assign mem[6641] = 5'h03;
  assign mem[6642] = 5'h12;
  assign mem[6643] = 5'h11;
  assign mem[6644] = 5'h10;
  assign mem[6645] = 5'h00;
  assign mem[6646] = 5'h01;
  assign mem[6647] = 5'h10;
  assign mem[6648] = 5'h00;
  assign mem[6649] = 5'h02;
  assign mem[6650] = 5'h11;
  assign mem[6651] = 5'h10;
  assign mem[6652] = 5'h00;
  assign mem[6653] = 5'h01;
  assign mem[6654] = 5'h10;
  assign mem[6655] = 5'h00;
  assign mem[6656] = 5'h08;
  assign mem[6657] = 5'h17;
  assign mem[6658] = 5'h16;
  assign mem[6659] = 5'h15;
  assign mem[6660] = 5'h14;
  assign mem[6661] = 5'h13;
  assign mem[6662] = 5'h12;
  assign mem[6663] = 5'h11;
  assign mem[6664] = 5'h10;
  assign mem[6665] = 5'h00;
  assign mem[6666] = 5'h01;
  assign mem[6667] = 5'h10;
  assign mem[6668] = 5'h00;
  assign mem[6669] = 5'h02;
  assign mem[6670] = 5'h11;
  assign mem[6671] = 5'h10;
  assign mem[6672] = 5'h00;
  assign mem[6673] = 5'h01;
  assign mem[6674] = 5'h10;
  assign mem[6675] = 5'h00;
  assign mem[6676] = 5'h03;
  assign mem[6677] = 5'h12;
  assign mem[6678] = 5'h11;
  assign mem[6679] = 5'h10;
  assign mem[6680] = 5'h00;
  assign mem[6681] = 5'h01;
  assign mem[6682] = 5'h10;
  assign mem[6683] = 5'h00;
  assign mem[6684] = 5'h02;
  assign mem[6685] = 5'h11;
  assign mem[6686] = 5'h10;
  assign mem[6687] = 5'h00;
  assign mem[6688] = 5'h01;
  assign mem[6689] = 5'h10;
  assign mem[6690] = 5'h00;
  assign mem[6691] = 5'h04;
  assign mem[6692] = 5'h13;
  assign mem[6693] = 5'h12;
  assign mem[6694] = 5'h11;
  assign mem[6695] = 5'h10;
  assign mem[6696] = 5'h00;
  assign mem[6697] = 5'h01;
  assign mem[6698] = 5'h10;
  assign mem[6699] = 5'h00;
  assign mem[6700] = 5'h02;
  assign mem[6701] = 5'h11;
  assign mem[6702] = 5'h10;
  assign mem[6703] = 5'h00;
  assign mem[6704] = 5'h01;
  assign mem[6705] = 5'h10;
  assign mem[6706] = 5'h00;
  assign mem[6707] = 5'h03;
  assign mem[6708] = 5'h12;
  assign mem[6709] = 5'h11;
  assign mem[6710] = 5'h10;
  assign mem[6711] = 5'h00;
  assign mem[6712] = 5'h01;
  assign mem[6713] = 5'h10;
  assign mem[6714] = 5'h00;
  assign mem[6715] = 5'h02;
  assign mem[6716] = 5'h11;
  assign mem[6717] = 5'h10;
  assign mem[6718] = 5'h00;
  assign mem[6719] = 5'h01;
  assign mem[6720] = 5'h10;
  assign mem[6721] = 5'h00;
  assign mem[6722] = 5'h05;
  assign mem[6723] = 5'h14;
  assign mem[6724] = 5'h13;
  assign mem[6725] = 5'h12;
  assign mem[6726] = 5'h11;
  assign mem[6727] = 5'h10;
  assign mem[6728] = 5'h00;
  assign mem[6729] = 5'h01;
  assign mem[6730] = 5'h10;
  assign mem[6731] = 5'h00;
  assign mem[6732] = 5'h02;
  assign mem[6733] = 5'h11;
  assign mem[6734] = 5'h10;
  assign mem[6735] = 5'h00;
  assign mem[6736] = 5'h01;
  assign mem[6737] = 5'h10;
  assign mem[6738] = 5'h00;
  assign mem[6739] = 5'h03;
  assign mem[6740] = 5'h12;
  assign mem[6741] = 5'h11;
  assign mem[6742] = 5'h10;
  assign mem[6743] = 5'h00;
  assign mem[6744] = 5'h01;
  assign mem[6745] = 5'h10;
  assign mem[6746] = 5'h00;
  assign mem[6747] = 5'h02;
  assign mem[6748] = 5'h11;
  assign mem[6749] = 5'h10;
  assign mem[6750] = 5'h00;
  assign mem[6751] = 5'h01;
  assign mem[6752] = 5'h10;
  assign mem[6753] = 5'h00;
  assign mem[6754] = 5'h04;
  assign mem[6755] = 5'h13;
  assign mem[6756] = 5'h12;
  assign mem[6757] = 5'h11;
  assign mem[6758] = 5'h10;
  assign mem[6759] = 5'h00;
  assign mem[6760] = 5'h01;
  assign mem[6761] = 5'h10;
  assign mem[6762] = 5'h00;
  assign mem[6763] = 5'h02;
  assign mem[6764] = 5'h11;
  assign mem[6765] = 5'h10;
  assign mem[6766] = 5'h00;
  assign mem[6767] = 5'h01;
  assign mem[6768] = 5'h10;
  assign mem[6769] = 5'h00;
  assign mem[6770] = 5'h03;
  assign mem[6771] = 5'h12;
  assign mem[6772] = 5'h11;
  assign mem[6773] = 5'h10;
  assign mem[6774] = 5'h00;
  assign mem[6775] = 5'h01;
  assign mem[6776] = 5'h10;
  assign mem[6777] = 5'h00;
  assign mem[6778] = 5'h02;
  assign mem[6779] = 5'h11;
  assign mem[6780] = 5'h10;
  assign mem[6781] = 5'h00;
  assign mem[6782] = 5'h01;
  assign mem[6783] = 5'h10;
  assign mem[6784] = 5'h00;
  assign mem[6785] = 5'h06;
  assign mem[6786] = 5'h15;
  assign mem[6787] = 5'h14;
  assign mem[6788] = 5'h13;
  assign mem[6789] = 5'h12;
  assign mem[6790] = 5'h11;
  assign mem[6791] = 5'h10;
  assign mem[6792] = 5'h00;
  assign mem[6793] = 5'h01;
  assign mem[6794] = 5'h10;
  assign mem[6795] = 5'h00;
  assign mem[6796] = 5'h02;
  assign mem[6797] = 5'h11;
  assign mem[6798] = 5'h10;
  assign mem[6799] = 5'h00;
  assign mem[6800] = 5'h01;
  assign mem[6801] = 5'h10;
  assign mem[6802] = 5'h00;
  assign mem[6803] = 5'h03;
  assign mem[6804] = 5'h12;
  assign mem[6805] = 5'h11;
  assign mem[6806] = 5'h10;
  assign mem[6807] = 5'h00;
  assign mem[6808] = 5'h01;
  assign mem[6809] = 5'h10;
  assign mem[6810] = 5'h00;
  assign mem[6811] = 5'h02;
  assign mem[6812] = 5'h11;
  assign mem[6813] = 5'h10;
  assign mem[6814] = 5'h00;
  assign mem[6815] = 5'h01;
  assign mem[6816] = 5'h10;
  assign mem[6817] = 5'h00;
  assign mem[6818] = 5'h04;
  assign mem[6819] = 5'h13;
  assign mem[6820] = 5'h12;
  assign mem[6821] = 5'h11;
  assign mem[6822] = 5'h10;
  assign mem[6823] = 5'h00;
  assign mem[6824] = 5'h01;
  assign mem[6825] = 5'h10;
  assign mem[6826] = 5'h00;
  assign mem[6827] = 5'h02;
  assign mem[6828] = 5'h11;
  assign mem[6829] = 5'h10;
  assign mem[6830] = 5'h00;
  assign mem[6831] = 5'h01;
  assign mem[6832] = 5'h10;
  assign mem[6833] = 5'h00;
  assign mem[6834] = 5'h03;
  assign mem[6835] = 5'h12;
  assign mem[6836] = 5'h11;
  assign mem[6837] = 5'h10;
  assign mem[6838] = 5'h00;
  assign mem[6839] = 5'h01;
  assign mem[6840] = 5'h10;
  assign mem[6841] = 5'h00;
  assign mem[6842] = 5'h02;
  assign mem[6843] = 5'h11;
  assign mem[6844] = 5'h10;
  assign mem[6845] = 5'h00;
  assign mem[6846] = 5'h01;
  assign mem[6847] = 5'h10;
  assign mem[6848] = 5'h00;
  assign mem[6849] = 5'h05;
  assign mem[6850] = 5'h14;
  assign mem[6851] = 5'h13;
  assign mem[6852] = 5'h12;
  assign mem[6853] = 5'h11;
  assign mem[6854] = 5'h10;
  assign mem[6855] = 5'h00;
  assign mem[6856] = 5'h01;
  assign mem[6857] = 5'h10;
  assign mem[6858] = 5'h00;
  assign mem[6859] = 5'h02;
  assign mem[6860] = 5'h11;
  assign mem[6861] = 5'h10;
  assign mem[6862] = 5'h00;
  assign mem[6863] = 5'h01;
  assign mem[6864] = 5'h10;
  assign mem[6865] = 5'h00;
  assign mem[6866] = 5'h03;
  assign mem[6867] = 5'h12;
  assign mem[6868] = 5'h11;
  assign mem[6869] = 5'h10;
  assign mem[6870] = 5'h00;
  assign mem[6871] = 5'h01;
  assign mem[6872] = 5'h10;
  assign mem[6873] = 5'h00;
  assign mem[6874] = 5'h02;
  assign mem[6875] = 5'h11;
  assign mem[6876] = 5'h10;
  assign mem[6877] = 5'h00;
  assign mem[6878] = 5'h01;
  assign mem[6879] = 5'h10;
  assign mem[6880] = 5'h00;
  assign mem[6881] = 5'h04;
  assign mem[6882] = 5'h13;
  assign mem[6883] = 5'h12;
  assign mem[6884] = 5'h11;
  assign mem[6885] = 5'h10;
  assign mem[6886] = 5'h00;
  assign mem[6887] = 5'h01;
  assign mem[6888] = 5'h10;
  assign mem[6889] = 5'h00;
  assign mem[6890] = 5'h02;
  assign mem[6891] = 5'h11;
  assign mem[6892] = 5'h10;
  assign mem[6893] = 5'h00;
  assign mem[6894] = 5'h01;
  assign mem[6895] = 5'h10;
  assign mem[6896] = 5'h00;
  assign mem[6897] = 5'h03;
  assign mem[6898] = 5'h12;
  assign mem[6899] = 5'h11;
  assign mem[6900] = 5'h10;
  assign mem[6901] = 5'h00;
  assign mem[6902] = 5'h01;
  assign mem[6903] = 5'h10;
  assign mem[6904] = 5'h00;
  assign mem[6905] = 5'h02;
  assign mem[6906] = 5'h11;
  assign mem[6907] = 5'h10;
  assign mem[6908] = 5'h00;
  assign mem[6909] = 5'h01;
  assign mem[6910] = 5'h10;
  assign mem[6911] = 5'h00;
  assign mem[6912] = 5'h07;
  assign mem[6913] = 5'h16;
  assign mem[6914] = 5'h15;
  assign mem[6915] = 5'h14;
  assign mem[6916] = 5'h13;
  assign mem[6917] = 5'h12;
  assign mem[6918] = 5'h11;
  assign mem[6919] = 5'h10;
  assign mem[6920] = 5'h00;
  assign mem[6921] = 5'h01;
  assign mem[6922] = 5'h10;
  assign mem[6923] = 5'h00;
  assign mem[6924] = 5'h02;
  assign mem[6925] = 5'h11;
  assign mem[6926] = 5'h10;
  assign mem[6927] = 5'h00;
  assign mem[6928] = 5'h01;
  assign mem[6929] = 5'h10;
  assign mem[6930] = 5'h00;
  assign mem[6931] = 5'h03;
  assign mem[6932] = 5'h12;
  assign mem[6933] = 5'h11;
  assign mem[6934] = 5'h10;
  assign mem[6935] = 5'h00;
  assign mem[6936] = 5'h01;
  assign mem[6937] = 5'h10;
  assign mem[6938] = 5'h00;
  assign mem[6939] = 5'h02;
  assign mem[6940] = 5'h11;
  assign mem[6941] = 5'h10;
  assign mem[6942] = 5'h00;
  assign mem[6943] = 5'h01;
  assign mem[6944] = 5'h10;
  assign mem[6945] = 5'h00;
  assign mem[6946] = 5'h04;
  assign mem[6947] = 5'h13;
  assign mem[6948] = 5'h12;
  assign mem[6949] = 5'h11;
  assign mem[6950] = 5'h10;
  assign mem[6951] = 5'h00;
  assign mem[6952] = 5'h01;
  assign mem[6953] = 5'h10;
  assign mem[6954] = 5'h00;
  assign mem[6955] = 5'h02;
  assign mem[6956] = 5'h11;
  assign mem[6957] = 5'h10;
  assign mem[6958] = 5'h00;
  assign mem[6959] = 5'h01;
  assign mem[6960] = 5'h10;
  assign mem[6961] = 5'h00;
  assign mem[6962] = 5'h03;
  assign mem[6963] = 5'h12;
  assign mem[6964] = 5'h11;
  assign mem[6965] = 5'h10;
  assign mem[6966] = 5'h00;
  assign mem[6967] = 5'h01;
  assign mem[6968] = 5'h10;
  assign mem[6969] = 5'h00;
  assign mem[6970] = 5'h02;
  assign mem[6971] = 5'h11;
  assign mem[6972] = 5'h10;
  assign mem[6973] = 5'h00;
  assign mem[6974] = 5'h01;
  assign mem[6975] = 5'h10;
  assign mem[6976] = 5'h00;
  assign mem[6977] = 5'h05;
  assign mem[6978] = 5'h14;
  assign mem[6979] = 5'h13;
  assign mem[6980] = 5'h12;
  assign mem[6981] = 5'h11;
  assign mem[6982] = 5'h10;
  assign mem[6983] = 5'h00;
  assign mem[6984] = 5'h01;
  assign mem[6985] = 5'h10;
  assign mem[6986] = 5'h00;
  assign mem[6987] = 5'h02;
  assign mem[6988] = 5'h11;
  assign mem[6989] = 5'h10;
  assign mem[6990] = 5'h00;
  assign mem[6991] = 5'h01;
  assign mem[6992] = 5'h10;
  assign mem[6993] = 5'h00;
  assign mem[6994] = 5'h03;
  assign mem[6995] = 5'h12;
  assign mem[6996] = 5'h11;
  assign mem[6997] = 5'h10;
  assign mem[6998] = 5'h00;
  assign mem[6999] = 5'h01;
  assign mem[7000] = 5'h10;
  assign mem[7001] = 5'h00;
  assign mem[7002] = 5'h02;
  assign mem[7003] = 5'h11;
  assign mem[7004] = 5'h10;
  assign mem[7005] = 5'h00;
  assign mem[7006] = 5'h01;
  assign mem[7007] = 5'h10;
  assign mem[7008] = 5'h00;
  assign mem[7009] = 5'h04;
  assign mem[7010] = 5'h13;
  assign mem[7011] = 5'h12;
  assign mem[7012] = 5'h11;
  assign mem[7013] = 5'h10;
  assign mem[7014] = 5'h00;
  assign mem[7015] = 5'h01;
  assign mem[7016] = 5'h10;
  assign mem[7017] = 5'h00;
  assign mem[7018] = 5'h02;
  assign mem[7019] = 5'h11;
  assign mem[7020] = 5'h10;
  assign mem[7021] = 5'h00;
  assign mem[7022] = 5'h01;
  assign mem[7023] = 5'h10;
  assign mem[7024] = 5'h00;
  assign mem[7025] = 5'h03;
  assign mem[7026] = 5'h12;
  assign mem[7027] = 5'h11;
  assign mem[7028] = 5'h10;
  assign mem[7029] = 5'h00;
  assign mem[7030] = 5'h01;
  assign mem[7031] = 5'h10;
  assign mem[7032] = 5'h00;
  assign mem[7033] = 5'h02;
  assign mem[7034] = 5'h11;
  assign mem[7035] = 5'h10;
  assign mem[7036] = 5'h00;
  assign mem[7037] = 5'h01;
  assign mem[7038] = 5'h10;
  assign mem[7039] = 5'h00;
  assign mem[7040] = 5'h06;
  assign mem[7041] = 5'h15;
  assign mem[7042] = 5'h14;
  assign mem[7043] = 5'h13;
  assign mem[7044] = 5'h12;
  assign mem[7045] = 5'h11;
  assign mem[7046] = 5'h10;
  assign mem[7047] = 5'h00;
  assign mem[7048] = 5'h01;
  assign mem[7049] = 5'h10;
  assign mem[7050] = 5'h00;
  assign mem[7051] = 5'h02;
  assign mem[7052] = 5'h11;
  assign mem[7053] = 5'h10;
  assign mem[7054] = 5'h00;
  assign mem[7055] = 5'h01;
  assign mem[7056] = 5'h10;
  assign mem[7057] = 5'h00;
  assign mem[7058] = 5'h03;
  assign mem[7059] = 5'h12;
  assign mem[7060] = 5'h11;
  assign mem[7061] = 5'h10;
  assign mem[7062] = 5'h00;
  assign mem[7063] = 5'h01;
  assign mem[7064] = 5'h10;
  assign mem[7065] = 5'h00;
  assign mem[7066] = 5'h02;
  assign mem[7067] = 5'h11;
  assign mem[7068] = 5'h10;
  assign mem[7069] = 5'h00;
  assign mem[7070] = 5'h01;
  assign mem[7071] = 5'h10;
  assign mem[7072] = 5'h00;
  assign mem[7073] = 5'h04;
  assign mem[7074] = 5'h13;
  assign mem[7075] = 5'h12;
  assign mem[7076] = 5'h11;
  assign mem[7077] = 5'h10;
  assign mem[7078] = 5'h00;
  assign mem[7079] = 5'h01;
  assign mem[7080] = 5'h10;
  assign mem[7081] = 5'h00;
  assign mem[7082] = 5'h02;
  assign mem[7083] = 5'h11;
  assign mem[7084] = 5'h10;
  assign mem[7085] = 5'h00;
  assign mem[7086] = 5'h01;
  assign mem[7087] = 5'h10;
  assign mem[7088] = 5'h00;
  assign mem[7089] = 5'h03;
  assign mem[7090] = 5'h12;
  assign mem[7091] = 5'h11;
  assign mem[7092] = 5'h10;
  assign mem[7093] = 5'h00;
  assign mem[7094] = 5'h01;
  assign mem[7095] = 5'h10;
  assign mem[7096] = 5'h00;
  assign mem[7097] = 5'h02;
  assign mem[7098] = 5'h11;
  assign mem[7099] = 5'h10;
  assign mem[7100] = 5'h00;
  assign mem[7101] = 5'h01;
  assign mem[7102] = 5'h10;
  assign mem[7103] = 5'h00;
  assign mem[7104] = 5'h05;
  assign mem[7105] = 5'h14;
  assign mem[7106] = 5'h13;
  assign mem[7107] = 5'h12;
  assign mem[7108] = 5'h11;
  assign mem[7109] = 5'h10;
  assign mem[7110] = 5'h00;
  assign mem[7111] = 5'h01;
  assign mem[7112] = 5'h10;
  assign mem[7113] = 5'h00;
  assign mem[7114] = 5'h02;
  assign mem[7115] = 5'h11;
  assign mem[7116] = 5'h10;
  assign mem[7117] = 5'h00;
  assign mem[7118] = 5'h01;
  assign mem[7119] = 5'h10;
  assign mem[7120] = 5'h00;
  assign mem[7121] = 5'h03;
  assign mem[7122] = 5'h12;
  assign mem[7123] = 5'h11;
  assign mem[7124] = 5'h10;
  assign mem[7125] = 5'h00;
  assign mem[7126] = 5'h01;
  assign mem[7127] = 5'h10;
  assign mem[7128] = 5'h00;
  assign mem[7129] = 5'h02;
  assign mem[7130] = 5'h11;
  assign mem[7131] = 5'h10;
  assign mem[7132] = 5'h00;
  assign mem[7133] = 5'h01;
  assign mem[7134] = 5'h10;
  assign mem[7135] = 5'h00;
  assign mem[7136] = 5'h04;
  assign mem[7137] = 5'h13;
  assign mem[7138] = 5'h12;
  assign mem[7139] = 5'h11;
  assign mem[7140] = 5'h10;
  assign mem[7141] = 5'h00;
  assign mem[7142] = 5'h01;
  assign mem[7143] = 5'h10;
  assign mem[7144] = 5'h00;
  assign mem[7145] = 5'h02;
  assign mem[7146] = 5'h11;
  assign mem[7147] = 5'h10;
  assign mem[7148] = 5'h00;
  assign mem[7149] = 5'h01;
  assign mem[7150] = 5'h10;
  assign mem[7151] = 5'h00;
  assign mem[7152] = 5'h03;
  assign mem[7153] = 5'h12;
  assign mem[7154] = 5'h11;
  assign mem[7155] = 5'h10;
  assign mem[7156] = 5'h00;
  assign mem[7157] = 5'h01;
  assign mem[7158] = 5'h10;
  assign mem[7159] = 5'h00;
  assign mem[7160] = 5'h02;
  assign mem[7161] = 5'h11;
  assign mem[7162] = 5'h10;
  assign mem[7163] = 5'h00;
  assign mem[7164] = 5'h01;
  assign mem[7165] = 5'h10;
  assign mem[7166] = 5'h00;
  assign mem[7167] = 5'h09;
  assign mem[7168] = 5'h18;
  assign mem[7169] = 5'h17;
  assign mem[7170] = 5'h16;
  assign mem[7171] = 5'h15;
  assign mem[7172] = 5'h14;
  assign mem[7173] = 5'h13;
  assign mem[7174] = 5'h12;
  assign mem[7175] = 5'h11;
  assign mem[7176] = 5'h10;
  assign mem[7177] = 5'h00;
  assign mem[7178] = 5'h01;
  assign mem[7179] = 5'h10;
  assign mem[7180] = 5'h00;
  assign mem[7181] = 5'h02;
  assign mem[7182] = 5'h11;
  assign mem[7183] = 5'h10;
  assign mem[7184] = 5'h00;
  assign mem[7185] = 5'h01;
  assign mem[7186] = 5'h10;
  assign mem[7187] = 5'h00;
  assign mem[7188] = 5'h03;
  assign mem[7189] = 5'h12;
  assign mem[7190] = 5'h11;
  assign mem[7191] = 5'h10;
  assign mem[7192] = 5'h00;
  assign mem[7193] = 5'h01;
  assign mem[7194] = 5'h10;
  assign mem[7195] = 5'h00;
  assign mem[7196] = 5'h02;
  assign mem[7197] = 5'h11;
  assign mem[7198] = 5'h10;
  assign mem[7199] = 5'h00;
  assign mem[7200] = 5'h01;
  assign mem[7201] = 5'h10;
  assign mem[7202] = 5'h00;
  assign mem[7203] = 5'h04;
  assign mem[7204] = 5'h13;
  assign mem[7205] = 5'h12;
  assign mem[7206] = 5'h11;
  assign mem[7207] = 5'h10;
  assign mem[7208] = 5'h00;
  assign mem[7209] = 5'h01;
  assign mem[7210] = 5'h10;
  assign mem[7211] = 5'h00;
  assign mem[7212] = 5'h02;
  assign mem[7213] = 5'h11;
  assign mem[7214] = 5'h10;
  assign mem[7215] = 5'h00;
  assign mem[7216] = 5'h01;
  assign mem[7217] = 5'h10;
  assign mem[7218] = 5'h00;
  assign mem[7219] = 5'h03;
  assign mem[7220] = 5'h12;
  assign mem[7221] = 5'h11;
  assign mem[7222] = 5'h10;
  assign mem[7223] = 5'h00;
  assign mem[7224] = 5'h01;
  assign mem[7225] = 5'h10;
  assign mem[7226] = 5'h00;
  assign mem[7227] = 5'h02;
  assign mem[7228] = 5'h11;
  assign mem[7229] = 5'h10;
  assign mem[7230] = 5'h00;
  assign mem[7231] = 5'h01;
  assign mem[7232] = 5'h10;
  assign mem[7233] = 5'h00;
  assign mem[7234] = 5'h05;
  assign mem[7235] = 5'h14;
  assign mem[7236] = 5'h13;
  assign mem[7237] = 5'h12;
  assign mem[7238] = 5'h11;
  assign mem[7239] = 5'h10;
  assign mem[7240] = 5'h00;
  assign mem[7241] = 5'h01;
  assign mem[7242] = 5'h10;
  assign mem[7243] = 5'h00;
  assign mem[7244] = 5'h02;
  assign mem[7245] = 5'h11;
  assign mem[7246] = 5'h10;
  assign mem[7247] = 5'h00;
  assign mem[7248] = 5'h01;
  assign mem[7249] = 5'h10;
  assign mem[7250] = 5'h00;
  assign mem[7251] = 5'h03;
  assign mem[7252] = 5'h12;
  assign mem[7253] = 5'h11;
  assign mem[7254] = 5'h10;
  assign mem[7255] = 5'h00;
  assign mem[7256] = 5'h01;
  assign mem[7257] = 5'h10;
  assign mem[7258] = 5'h00;
  assign mem[7259] = 5'h02;
  assign mem[7260] = 5'h11;
  assign mem[7261] = 5'h10;
  assign mem[7262] = 5'h00;
  assign mem[7263] = 5'h01;
  assign mem[7264] = 5'h10;
  assign mem[7265] = 5'h00;
  assign mem[7266] = 5'h04;
  assign mem[7267] = 5'h13;
  assign mem[7268] = 5'h12;
  assign mem[7269] = 5'h11;
  assign mem[7270] = 5'h10;
  assign mem[7271] = 5'h00;
  assign mem[7272] = 5'h01;
  assign mem[7273] = 5'h10;
  assign mem[7274] = 5'h00;
  assign mem[7275] = 5'h02;
  assign mem[7276] = 5'h11;
  assign mem[7277] = 5'h10;
  assign mem[7278] = 5'h00;
  assign mem[7279] = 5'h01;
  assign mem[7280] = 5'h10;
  assign mem[7281] = 5'h00;
  assign mem[7282] = 5'h03;
  assign mem[7283] = 5'h12;
  assign mem[7284] = 5'h11;
  assign mem[7285] = 5'h10;
  assign mem[7286] = 5'h00;
  assign mem[7287] = 5'h01;
  assign mem[7288] = 5'h10;
  assign mem[7289] = 5'h00;
  assign mem[7290] = 5'h02;
  assign mem[7291] = 5'h11;
  assign mem[7292] = 5'h10;
  assign mem[7293] = 5'h00;
  assign mem[7294] = 5'h01;
  assign mem[7295] = 5'h10;
  assign mem[7296] = 5'h00;
  assign mem[7297] = 5'h06;
  assign mem[7298] = 5'h15;
  assign mem[7299] = 5'h14;
  assign mem[7300] = 5'h13;
  assign mem[7301] = 5'h12;
  assign mem[7302] = 5'h11;
  assign mem[7303] = 5'h10;
  assign mem[7304] = 5'h00;
  assign mem[7305] = 5'h01;
  assign mem[7306] = 5'h10;
  assign mem[7307] = 5'h00;
  assign mem[7308] = 5'h02;
  assign mem[7309] = 5'h11;
  assign mem[7310] = 5'h10;
  assign mem[7311] = 5'h00;
  assign mem[7312] = 5'h01;
  assign mem[7313] = 5'h10;
  assign mem[7314] = 5'h00;
  assign mem[7315] = 5'h03;
  assign mem[7316] = 5'h12;
  assign mem[7317] = 5'h11;
  assign mem[7318] = 5'h10;
  assign mem[7319] = 5'h00;
  assign mem[7320] = 5'h01;
  assign mem[7321] = 5'h10;
  assign mem[7322] = 5'h00;
  assign mem[7323] = 5'h02;
  assign mem[7324] = 5'h11;
  assign mem[7325] = 5'h10;
  assign mem[7326] = 5'h00;
  assign mem[7327] = 5'h01;
  assign mem[7328] = 5'h10;
  assign mem[7329] = 5'h00;
  assign mem[7330] = 5'h04;
  assign mem[7331] = 5'h13;
  assign mem[7332] = 5'h12;
  assign mem[7333] = 5'h11;
  assign mem[7334] = 5'h10;
  assign mem[7335] = 5'h00;
  assign mem[7336] = 5'h01;
  assign mem[7337] = 5'h10;
  assign mem[7338] = 5'h00;
  assign mem[7339] = 5'h02;
  assign mem[7340] = 5'h11;
  assign mem[7341] = 5'h10;
  assign mem[7342] = 5'h00;
  assign mem[7343] = 5'h01;
  assign mem[7344] = 5'h10;
  assign mem[7345] = 5'h00;
  assign mem[7346] = 5'h03;
  assign mem[7347] = 5'h12;
  assign mem[7348] = 5'h11;
  assign mem[7349] = 5'h10;
  assign mem[7350] = 5'h00;
  assign mem[7351] = 5'h01;
  assign mem[7352] = 5'h10;
  assign mem[7353] = 5'h00;
  assign mem[7354] = 5'h02;
  assign mem[7355] = 5'h11;
  assign mem[7356] = 5'h10;
  assign mem[7357] = 5'h00;
  assign mem[7358] = 5'h01;
  assign mem[7359] = 5'h10;
  assign mem[7360] = 5'h00;
  assign mem[7361] = 5'h05;
  assign mem[7362] = 5'h14;
  assign mem[7363] = 5'h13;
  assign mem[7364] = 5'h12;
  assign mem[7365] = 5'h11;
  assign mem[7366] = 5'h10;
  assign mem[7367] = 5'h00;
  assign mem[7368] = 5'h01;
  assign mem[7369] = 5'h10;
  assign mem[7370] = 5'h00;
  assign mem[7371] = 5'h02;
  assign mem[7372] = 5'h11;
  assign mem[7373] = 5'h10;
  assign mem[7374] = 5'h00;
  assign mem[7375] = 5'h01;
  assign mem[7376] = 5'h10;
  assign mem[7377] = 5'h00;
  assign mem[7378] = 5'h03;
  assign mem[7379] = 5'h12;
  assign mem[7380] = 5'h11;
  assign mem[7381] = 5'h10;
  assign mem[7382] = 5'h00;
  assign mem[7383] = 5'h01;
  assign mem[7384] = 5'h10;
  assign mem[7385] = 5'h00;
  assign mem[7386] = 5'h02;
  assign mem[7387] = 5'h11;
  assign mem[7388] = 5'h10;
  assign mem[7389] = 5'h00;
  assign mem[7390] = 5'h01;
  assign mem[7391] = 5'h10;
  assign mem[7392] = 5'h00;
  assign mem[7393] = 5'h04;
  assign mem[7394] = 5'h13;
  assign mem[7395] = 5'h12;
  assign mem[7396] = 5'h11;
  assign mem[7397] = 5'h10;
  assign mem[7398] = 5'h00;
  assign mem[7399] = 5'h01;
  assign mem[7400] = 5'h10;
  assign mem[7401] = 5'h00;
  assign mem[7402] = 5'h02;
  assign mem[7403] = 5'h11;
  assign mem[7404] = 5'h10;
  assign mem[7405] = 5'h00;
  assign mem[7406] = 5'h01;
  assign mem[7407] = 5'h10;
  assign mem[7408] = 5'h00;
  assign mem[7409] = 5'h03;
  assign mem[7410] = 5'h12;
  assign mem[7411] = 5'h11;
  assign mem[7412] = 5'h10;
  assign mem[7413] = 5'h00;
  assign mem[7414] = 5'h01;
  assign mem[7415] = 5'h10;
  assign mem[7416] = 5'h00;
  assign mem[7417] = 5'h02;
  assign mem[7418] = 5'h11;
  assign mem[7419] = 5'h10;
  assign mem[7420] = 5'h00;
  assign mem[7421] = 5'h01;
  assign mem[7422] = 5'h10;
  assign mem[7423] = 5'h00;
  assign mem[7424] = 5'h07;
  assign mem[7425] = 5'h16;
  assign mem[7426] = 5'h15;
  assign mem[7427] = 5'h14;
  assign mem[7428] = 5'h13;
  assign mem[7429] = 5'h12;
  assign mem[7430] = 5'h11;
  assign mem[7431] = 5'h10;
  assign mem[7432] = 5'h00;
  assign mem[7433] = 5'h01;
  assign mem[7434] = 5'h10;
  assign mem[7435] = 5'h00;
  assign mem[7436] = 5'h02;
  assign mem[7437] = 5'h11;
  assign mem[7438] = 5'h10;
  assign mem[7439] = 5'h00;
  assign mem[7440] = 5'h01;
  assign mem[7441] = 5'h10;
  assign mem[7442] = 5'h00;
  assign mem[7443] = 5'h03;
  assign mem[7444] = 5'h12;
  assign mem[7445] = 5'h11;
  assign mem[7446] = 5'h10;
  assign mem[7447] = 5'h00;
  assign mem[7448] = 5'h01;
  assign mem[7449] = 5'h10;
  assign mem[7450] = 5'h00;
  assign mem[7451] = 5'h02;
  assign mem[7452] = 5'h11;
  assign mem[7453] = 5'h10;
  assign mem[7454] = 5'h00;
  assign mem[7455] = 5'h01;
  assign mem[7456] = 5'h10;
  assign mem[7457] = 5'h00;
  assign mem[7458] = 5'h04;
  assign mem[7459] = 5'h13;
  assign mem[7460] = 5'h12;
  assign mem[7461] = 5'h11;
  assign mem[7462] = 5'h10;
  assign mem[7463] = 5'h00;
  assign mem[7464] = 5'h01;
  assign mem[7465] = 5'h10;
  assign mem[7466] = 5'h00;
  assign mem[7467] = 5'h02;
  assign mem[7468] = 5'h11;
  assign mem[7469] = 5'h10;
  assign mem[7470] = 5'h00;
  assign mem[7471] = 5'h01;
  assign mem[7472] = 5'h10;
  assign mem[7473] = 5'h00;
  assign mem[7474] = 5'h03;
  assign mem[7475] = 5'h12;
  assign mem[7476] = 5'h11;
  assign mem[7477] = 5'h10;
  assign mem[7478] = 5'h00;
  assign mem[7479] = 5'h01;
  assign mem[7480] = 5'h10;
  assign mem[7481] = 5'h00;
  assign mem[7482] = 5'h02;
  assign mem[7483] = 5'h11;
  assign mem[7484] = 5'h10;
  assign mem[7485] = 5'h00;
  assign mem[7486] = 5'h01;
  assign mem[7487] = 5'h10;
  assign mem[7488] = 5'h00;
  assign mem[7489] = 5'h05;
  assign mem[7490] = 5'h14;
  assign mem[7491] = 5'h13;
  assign mem[7492] = 5'h12;
  assign mem[7493] = 5'h11;
  assign mem[7494] = 5'h10;
  assign mem[7495] = 5'h00;
  assign mem[7496] = 5'h01;
  assign mem[7497] = 5'h10;
  assign mem[7498] = 5'h00;
  assign mem[7499] = 5'h02;
  assign mem[7500] = 5'h11;
  assign mem[7501] = 5'h10;
  assign mem[7502] = 5'h00;
  assign mem[7503] = 5'h01;
  assign mem[7504] = 5'h10;
  assign mem[7505] = 5'h00;
  assign mem[7506] = 5'h03;
  assign mem[7507] = 5'h12;
  assign mem[7508] = 5'h11;
  assign mem[7509] = 5'h10;
  assign mem[7510] = 5'h00;
  assign mem[7511] = 5'h01;
  assign mem[7512] = 5'h10;
  assign mem[7513] = 5'h00;
  assign mem[7514] = 5'h02;
  assign mem[7515] = 5'h11;
  assign mem[7516] = 5'h10;
  assign mem[7517] = 5'h00;
  assign mem[7518] = 5'h01;
  assign mem[7519] = 5'h10;
  assign mem[7520] = 5'h00;
  assign mem[7521] = 5'h04;
  assign mem[7522] = 5'h13;
  assign mem[7523] = 5'h12;
  assign mem[7524] = 5'h11;
  assign mem[7525] = 5'h10;
  assign mem[7526] = 5'h00;
  assign mem[7527] = 5'h01;
  assign mem[7528] = 5'h10;
  assign mem[7529] = 5'h00;
  assign mem[7530] = 5'h02;
  assign mem[7531] = 5'h11;
  assign mem[7532] = 5'h10;
  assign mem[7533] = 5'h00;
  assign mem[7534] = 5'h01;
  assign mem[7535] = 5'h10;
  assign mem[7536] = 5'h00;
  assign mem[7537] = 5'h03;
  assign mem[7538] = 5'h12;
  assign mem[7539] = 5'h11;
  assign mem[7540] = 5'h10;
  assign mem[7541] = 5'h00;
  assign mem[7542] = 5'h01;
  assign mem[7543] = 5'h10;
  assign mem[7544] = 5'h00;
  assign mem[7545] = 5'h02;
  assign mem[7546] = 5'h11;
  assign mem[7547] = 5'h10;
  assign mem[7548] = 5'h00;
  assign mem[7549] = 5'h01;
  assign mem[7550] = 5'h10;
  assign mem[7551] = 5'h00;
  assign mem[7552] = 5'h06;
  assign mem[7553] = 5'h15;
  assign mem[7554] = 5'h14;
  assign mem[7555] = 5'h13;
  assign mem[7556] = 5'h12;
  assign mem[7557] = 5'h11;
  assign mem[7558] = 5'h10;
  assign mem[7559] = 5'h00;
  assign mem[7560] = 5'h01;
  assign mem[7561] = 5'h10;
  assign mem[7562] = 5'h00;
  assign mem[7563] = 5'h02;
  assign mem[7564] = 5'h11;
  assign mem[7565] = 5'h10;
  assign mem[7566] = 5'h00;
  assign mem[7567] = 5'h01;
  assign mem[7568] = 5'h10;
  assign mem[7569] = 5'h00;
  assign mem[7570] = 5'h03;
  assign mem[7571] = 5'h12;
  assign mem[7572] = 5'h11;
  assign mem[7573] = 5'h10;
  assign mem[7574] = 5'h00;
  assign mem[7575] = 5'h01;
  assign mem[7576] = 5'h10;
  assign mem[7577] = 5'h00;
  assign mem[7578] = 5'h02;
  assign mem[7579] = 5'h11;
  assign mem[7580] = 5'h10;
  assign mem[7581] = 5'h00;
  assign mem[7582] = 5'h01;
  assign mem[7583] = 5'h10;
  assign mem[7584] = 5'h00;
  assign mem[7585] = 5'h04;
  assign mem[7586] = 5'h13;
  assign mem[7587] = 5'h12;
  assign mem[7588] = 5'h11;
  assign mem[7589] = 5'h10;
  assign mem[7590] = 5'h00;
  assign mem[7591] = 5'h01;
  assign mem[7592] = 5'h10;
  assign mem[7593] = 5'h00;
  assign mem[7594] = 5'h02;
  assign mem[7595] = 5'h11;
  assign mem[7596] = 5'h10;
  assign mem[7597] = 5'h00;
  assign mem[7598] = 5'h01;
  assign mem[7599] = 5'h10;
  assign mem[7600] = 5'h00;
  assign mem[7601] = 5'h03;
  assign mem[7602] = 5'h12;
  assign mem[7603] = 5'h11;
  assign mem[7604] = 5'h10;
  assign mem[7605] = 5'h00;
  assign mem[7606] = 5'h01;
  assign mem[7607] = 5'h10;
  assign mem[7608] = 5'h00;
  assign mem[7609] = 5'h02;
  assign mem[7610] = 5'h11;
  assign mem[7611] = 5'h10;
  assign mem[7612] = 5'h00;
  assign mem[7613] = 5'h01;
  assign mem[7614] = 5'h10;
  assign mem[7615] = 5'h00;
  assign mem[7616] = 5'h05;
  assign mem[7617] = 5'h14;
  assign mem[7618] = 5'h13;
  assign mem[7619] = 5'h12;
  assign mem[7620] = 5'h11;
  assign mem[7621] = 5'h10;
  assign mem[7622] = 5'h00;
  assign mem[7623] = 5'h01;
  assign mem[7624] = 5'h10;
  assign mem[7625] = 5'h00;
  assign mem[7626] = 5'h02;
  assign mem[7627] = 5'h11;
  assign mem[7628] = 5'h10;
  assign mem[7629] = 5'h00;
  assign mem[7630] = 5'h01;
  assign mem[7631] = 5'h10;
  assign mem[7632] = 5'h00;
  assign mem[7633] = 5'h03;
  assign mem[7634] = 5'h12;
  assign mem[7635] = 5'h11;
  assign mem[7636] = 5'h10;
  assign mem[7637] = 5'h00;
  assign mem[7638] = 5'h01;
  assign mem[7639] = 5'h10;
  assign mem[7640] = 5'h00;
  assign mem[7641] = 5'h02;
  assign mem[7642] = 5'h11;
  assign mem[7643] = 5'h10;
  assign mem[7644] = 5'h00;
  assign mem[7645] = 5'h01;
  assign mem[7646] = 5'h10;
  assign mem[7647] = 5'h00;
  assign mem[7648] = 5'h04;
  assign mem[7649] = 5'h13;
  assign mem[7650] = 5'h12;
  assign mem[7651] = 5'h11;
  assign mem[7652] = 5'h10;
  assign mem[7653] = 5'h00;
  assign mem[7654] = 5'h01;
  assign mem[7655] = 5'h10;
  assign mem[7656] = 5'h00;
  assign mem[7657] = 5'h02;
  assign mem[7658] = 5'h11;
  assign mem[7659] = 5'h10;
  assign mem[7660] = 5'h00;
  assign mem[7661] = 5'h01;
  assign mem[7662] = 5'h10;
  assign mem[7663] = 5'h00;
  assign mem[7664] = 5'h03;
  assign mem[7665] = 5'h12;
  assign mem[7666] = 5'h11;
  assign mem[7667] = 5'h10;
  assign mem[7668] = 5'h00;
  assign mem[7669] = 5'h01;
  assign mem[7670] = 5'h10;
  assign mem[7671] = 5'h00;
  assign mem[7672] = 5'h02;
  assign mem[7673] = 5'h11;
  assign mem[7674] = 5'h10;
  assign mem[7675] = 5'h00;
  assign mem[7676] = 5'h01;
  assign mem[7677] = 5'h10;
  assign mem[7678] = 5'h00;
  assign mem[7679] = 5'h08;
  assign mem[7680] = 5'h17;
  assign mem[7681] = 5'h16;
  assign mem[7682] = 5'h15;
  assign mem[7683] = 5'h14;
  assign mem[7684] = 5'h13;
  assign mem[7685] = 5'h12;
  assign mem[7686] = 5'h11;
  assign mem[7687] = 5'h10;
  assign mem[7688] = 5'h00;
  assign mem[7689] = 5'h01;
  assign mem[7690] = 5'h10;
  assign mem[7691] = 5'h00;
  assign mem[7692] = 5'h02;
  assign mem[7693] = 5'h11;
  assign mem[7694] = 5'h10;
  assign mem[7695] = 5'h00;
  assign mem[7696] = 5'h01;
  assign mem[7697] = 5'h10;
  assign mem[7698] = 5'h00;
  assign mem[7699] = 5'h03;
  assign mem[7700] = 5'h12;
  assign mem[7701] = 5'h11;
  assign mem[7702] = 5'h10;
  assign mem[7703] = 5'h00;
  assign mem[7704] = 5'h01;
  assign mem[7705] = 5'h10;
  assign mem[7706] = 5'h00;
  assign mem[7707] = 5'h02;
  assign mem[7708] = 5'h11;
  assign mem[7709] = 5'h10;
  assign mem[7710] = 5'h00;
  assign mem[7711] = 5'h01;
  assign mem[7712] = 5'h10;
  assign mem[7713] = 5'h00;
  assign mem[7714] = 5'h04;
  assign mem[7715] = 5'h13;
  assign mem[7716] = 5'h12;
  assign mem[7717] = 5'h11;
  assign mem[7718] = 5'h10;
  assign mem[7719] = 5'h00;
  assign mem[7720] = 5'h01;
  assign mem[7721] = 5'h10;
  assign mem[7722] = 5'h00;
  assign mem[7723] = 5'h02;
  assign mem[7724] = 5'h11;
  assign mem[7725] = 5'h10;
  assign mem[7726] = 5'h00;
  assign mem[7727] = 5'h01;
  assign mem[7728] = 5'h10;
  assign mem[7729] = 5'h00;
  assign mem[7730] = 5'h03;
  assign mem[7731] = 5'h12;
  assign mem[7732] = 5'h11;
  assign mem[7733] = 5'h10;
  assign mem[7734] = 5'h00;
  assign mem[7735] = 5'h01;
  assign mem[7736] = 5'h10;
  assign mem[7737] = 5'h00;
  assign mem[7738] = 5'h02;
  assign mem[7739] = 5'h11;
  assign mem[7740] = 5'h10;
  assign mem[7741] = 5'h00;
  assign mem[7742] = 5'h01;
  assign mem[7743] = 5'h10;
  assign mem[7744] = 5'h00;
  assign mem[7745] = 5'h05;
  assign mem[7746] = 5'h14;
  assign mem[7747] = 5'h13;
  assign mem[7748] = 5'h12;
  assign mem[7749] = 5'h11;
  assign mem[7750] = 5'h10;
  assign mem[7751] = 5'h00;
  assign mem[7752] = 5'h01;
  assign mem[7753] = 5'h10;
  assign mem[7754] = 5'h00;
  assign mem[7755] = 5'h02;
  assign mem[7756] = 5'h11;
  assign mem[7757] = 5'h10;
  assign mem[7758] = 5'h00;
  assign mem[7759] = 5'h01;
  assign mem[7760] = 5'h10;
  assign mem[7761] = 5'h00;
  assign mem[7762] = 5'h03;
  assign mem[7763] = 5'h12;
  assign mem[7764] = 5'h11;
  assign mem[7765] = 5'h10;
  assign mem[7766] = 5'h00;
  assign mem[7767] = 5'h01;
  assign mem[7768] = 5'h10;
  assign mem[7769] = 5'h00;
  assign mem[7770] = 5'h02;
  assign mem[7771] = 5'h11;
  assign mem[7772] = 5'h10;
  assign mem[7773] = 5'h00;
  assign mem[7774] = 5'h01;
  assign mem[7775] = 5'h10;
  assign mem[7776] = 5'h00;
  assign mem[7777] = 5'h04;
  assign mem[7778] = 5'h13;
  assign mem[7779] = 5'h12;
  assign mem[7780] = 5'h11;
  assign mem[7781] = 5'h10;
  assign mem[7782] = 5'h00;
  assign mem[7783] = 5'h01;
  assign mem[7784] = 5'h10;
  assign mem[7785] = 5'h00;
  assign mem[7786] = 5'h02;
  assign mem[7787] = 5'h11;
  assign mem[7788] = 5'h10;
  assign mem[7789] = 5'h00;
  assign mem[7790] = 5'h01;
  assign mem[7791] = 5'h10;
  assign mem[7792] = 5'h00;
  assign mem[7793] = 5'h03;
  assign mem[7794] = 5'h12;
  assign mem[7795] = 5'h11;
  assign mem[7796] = 5'h10;
  assign mem[7797] = 5'h00;
  assign mem[7798] = 5'h01;
  assign mem[7799] = 5'h10;
  assign mem[7800] = 5'h00;
  assign mem[7801] = 5'h02;
  assign mem[7802] = 5'h11;
  assign mem[7803] = 5'h10;
  assign mem[7804] = 5'h00;
  assign mem[7805] = 5'h01;
  assign mem[7806] = 5'h10;
  assign mem[7807] = 5'h00;
  assign mem[7808] = 5'h06;
  assign mem[7809] = 5'h15;
  assign mem[7810] = 5'h14;
  assign mem[7811] = 5'h13;
  assign mem[7812] = 5'h12;
  assign mem[7813] = 5'h11;
  assign mem[7814] = 5'h10;
  assign mem[7815] = 5'h00;
  assign mem[7816] = 5'h01;
  assign mem[7817] = 5'h10;
  assign mem[7818] = 5'h00;
  assign mem[7819] = 5'h02;
  assign mem[7820] = 5'h11;
  assign mem[7821] = 5'h10;
  assign mem[7822] = 5'h00;
  assign mem[7823] = 5'h01;
  assign mem[7824] = 5'h10;
  assign mem[7825] = 5'h00;
  assign mem[7826] = 5'h03;
  assign mem[7827] = 5'h12;
  assign mem[7828] = 5'h11;
  assign mem[7829] = 5'h10;
  assign mem[7830] = 5'h00;
  assign mem[7831] = 5'h01;
  assign mem[7832] = 5'h10;
  assign mem[7833] = 5'h00;
  assign mem[7834] = 5'h02;
  assign mem[7835] = 5'h11;
  assign mem[7836] = 5'h10;
  assign mem[7837] = 5'h00;
  assign mem[7838] = 5'h01;
  assign mem[7839] = 5'h10;
  assign mem[7840] = 5'h00;
  assign mem[7841] = 5'h04;
  assign mem[7842] = 5'h13;
  assign mem[7843] = 5'h12;
  assign mem[7844] = 5'h11;
  assign mem[7845] = 5'h10;
  assign mem[7846] = 5'h00;
  assign mem[7847] = 5'h01;
  assign mem[7848] = 5'h10;
  assign mem[7849] = 5'h00;
  assign mem[7850] = 5'h02;
  assign mem[7851] = 5'h11;
  assign mem[7852] = 5'h10;
  assign mem[7853] = 5'h00;
  assign mem[7854] = 5'h01;
  assign mem[7855] = 5'h10;
  assign mem[7856] = 5'h00;
  assign mem[7857] = 5'h03;
  assign mem[7858] = 5'h12;
  assign mem[7859] = 5'h11;
  assign mem[7860] = 5'h10;
  assign mem[7861] = 5'h00;
  assign mem[7862] = 5'h01;
  assign mem[7863] = 5'h10;
  assign mem[7864] = 5'h00;
  assign mem[7865] = 5'h02;
  assign mem[7866] = 5'h11;
  assign mem[7867] = 5'h10;
  assign mem[7868] = 5'h00;
  assign mem[7869] = 5'h01;
  assign mem[7870] = 5'h10;
  assign mem[7871] = 5'h00;
  assign mem[7872] = 5'h05;
  assign mem[7873] = 5'h14;
  assign mem[7874] = 5'h13;
  assign mem[7875] = 5'h12;
  assign mem[7876] = 5'h11;
  assign mem[7877] = 5'h10;
  assign mem[7878] = 5'h00;
  assign mem[7879] = 5'h01;
  assign mem[7880] = 5'h10;
  assign mem[7881] = 5'h00;
  assign mem[7882] = 5'h02;
  assign mem[7883] = 5'h11;
  assign mem[7884] = 5'h10;
  assign mem[7885] = 5'h00;
  assign mem[7886] = 5'h01;
  assign mem[7887] = 5'h10;
  assign mem[7888] = 5'h00;
  assign mem[7889] = 5'h03;
  assign mem[7890] = 5'h12;
  assign mem[7891] = 5'h11;
  assign mem[7892] = 5'h10;
  assign mem[7893] = 5'h00;
  assign mem[7894] = 5'h01;
  assign mem[7895] = 5'h10;
  assign mem[7896] = 5'h00;
  assign mem[7897] = 5'h02;
  assign mem[7898] = 5'h11;
  assign mem[7899] = 5'h10;
  assign mem[7900] = 5'h00;
  assign mem[7901] = 5'h01;
  assign mem[7902] = 5'h10;
  assign mem[7903] = 5'h00;
  assign mem[7904] = 5'h04;
  assign mem[7905] = 5'h13;
  assign mem[7906] = 5'h12;
  assign mem[7907] = 5'h11;
  assign mem[7908] = 5'h10;
  assign mem[7909] = 5'h00;
  assign mem[7910] = 5'h01;
  assign mem[7911] = 5'h10;
  assign mem[7912] = 5'h00;
  assign mem[7913] = 5'h02;
  assign mem[7914] = 5'h11;
  assign mem[7915] = 5'h10;
  assign mem[7916] = 5'h00;
  assign mem[7917] = 5'h01;
  assign mem[7918] = 5'h10;
  assign mem[7919] = 5'h00;
  assign mem[7920] = 5'h03;
  assign mem[7921] = 5'h12;
  assign mem[7922] = 5'h11;
  assign mem[7923] = 5'h10;
  assign mem[7924] = 5'h00;
  assign mem[7925] = 5'h01;
  assign mem[7926] = 5'h10;
  assign mem[7927] = 5'h00;
  assign mem[7928] = 5'h02;
  assign mem[7929] = 5'h11;
  assign mem[7930] = 5'h10;
  assign mem[7931] = 5'h00;
  assign mem[7932] = 5'h01;
  assign mem[7933] = 5'h10;
  assign mem[7934] = 5'h00;
  assign mem[7935] = 5'h07;
  assign mem[7936] = 5'h16;
  assign mem[7937] = 5'h15;
  assign mem[7938] = 5'h14;
  assign mem[7939] = 5'h13;
  assign mem[7940] = 5'h12;
  assign mem[7941] = 5'h11;
  assign mem[7942] = 5'h10;
  assign mem[7943] = 5'h00;
  assign mem[7944] = 5'h01;
  assign mem[7945] = 5'h10;
  assign mem[7946] = 5'h00;
  assign mem[7947] = 5'h02;
  assign mem[7948] = 5'h11;
  assign mem[7949] = 5'h10;
  assign mem[7950] = 5'h00;
  assign mem[7951] = 5'h01;
  assign mem[7952] = 5'h10;
  assign mem[7953] = 5'h00;
  assign mem[7954] = 5'h03;
  assign mem[7955] = 5'h12;
  assign mem[7956] = 5'h11;
  assign mem[7957] = 5'h10;
  assign mem[7958] = 5'h00;
  assign mem[7959] = 5'h01;
  assign mem[7960] = 5'h10;
  assign mem[7961] = 5'h00;
  assign mem[7962] = 5'h02;
  assign mem[7963] = 5'h11;
  assign mem[7964] = 5'h10;
  assign mem[7965] = 5'h00;
  assign mem[7966] = 5'h01;
  assign mem[7967] = 5'h10;
  assign mem[7968] = 5'h00;
  assign mem[7969] = 5'h04;
  assign mem[7970] = 5'h13;
  assign mem[7971] = 5'h12;
  assign mem[7972] = 5'h11;
  assign mem[7973] = 5'h10;
  assign mem[7974] = 5'h00;
  assign mem[7975] = 5'h01;
  assign mem[7976] = 5'h10;
  assign mem[7977] = 5'h00;
  assign mem[7978] = 5'h02;
  assign mem[7979] = 5'h11;
  assign mem[7980] = 5'h10;
  assign mem[7981] = 5'h00;
  assign mem[7982] = 5'h01;
  assign mem[7983] = 5'h10;
  assign mem[7984] = 5'h00;
  assign mem[7985] = 5'h03;
  assign mem[7986] = 5'h12;
  assign mem[7987] = 5'h11;
  assign mem[7988] = 5'h10;
  assign mem[7989] = 5'h00;
  assign mem[7990] = 5'h01;
  assign mem[7991] = 5'h10;
  assign mem[7992] = 5'h00;
  assign mem[7993] = 5'h02;
  assign mem[7994] = 5'h11;
  assign mem[7995] = 5'h10;
  assign mem[7996] = 5'h00;
  assign mem[7997] = 5'h01;
  assign mem[7998] = 5'h10;
  assign mem[7999] = 5'h00;
  assign mem[8000] = 5'h05;
  assign mem[8001] = 5'h14;
  assign mem[8002] = 5'h13;
  assign mem[8003] = 5'h12;
  assign mem[8004] = 5'h11;
  assign mem[8005] = 5'h10;
  assign mem[8006] = 5'h00;
  assign mem[8007] = 5'h01;
  assign mem[8008] = 5'h10;
  assign mem[8009] = 5'h00;
  assign mem[8010] = 5'h02;
  assign mem[8011] = 5'h11;
  assign mem[8012] = 5'h10;
  assign mem[8013] = 5'h00;
  assign mem[8014] = 5'h01;
  assign mem[8015] = 5'h10;
  assign mem[8016] = 5'h00;
  assign mem[8017] = 5'h03;
  assign mem[8018] = 5'h12;
  assign mem[8019] = 5'h11;
  assign mem[8020] = 5'h10;
  assign mem[8021] = 5'h00;
  assign mem[8022] = 5'h01;
  assign mem[8023] = 5'h10;
  assign mem[8024] = 5'h00;
  assign mem[8025] = 5'h02;
  assign mem[8026] = 5'h11;
  assign mem[8027] = 5'h10;
  assign mem[8028] = 5'h00;
  assign mem[8029] = 5'h01;
  assign mem[8030] = 5'h10;
  assign mem[8031] = 5'h00;
  assign mem[8032] = 5'h04;
  assign mem[8033] = 5'h13;
  assign mem[8034] = 5'h12;
  assign mem[8035] = 5'h11;
  assign mem[8036] = 5'h10;
  assign mem[8037] = 5'h00;
  assign mem[8038] = 5'h01;
  assign mem[8039] = 5'h10;
  assign mem[8040] = 5'h00;
  assign mem[8041] = 5'h02;
  assign mem[8042] = 5'h11;
  assign mem[8043] = 5'h10;
  assign mem[8044] = 5'h00;
  assign mem[8045] = 5'h01;
  assign mem[8046] = 5'h10;
  assign mem[8047] = 5'h00;
  assign mem[8048] = 5'h03;
  assign mem[8049] = 5'h12;
  assign mem[8050] = 5'h11;
  assign mem[8051] = 5'h10;
  assign mem[8052] = 5'h00;
  assign mem[8053] = 5'h01;
  assign mem[8054] = 5'h10;
  assign mem[8055] = 5'h00;
  assign mem[8056] = 5'h02;
  assign mem[8057] = 5'h11;
  assign mem[8058] = 5'h10;
  assign mem[8059] = 5'h00;
  assign mem[8060] = 5'h01;
  assign mem[8061] = 5'h10;
  assign mem[8062] = 5'h00;
  assign mem[8063] = 5'h06;
  assign mem[8064] = 5'h15;
  assign mem[8065] = 5'h14;
  assign mem[8066] = 5'h13;
  assign mem[8067] = 5'h12;
  assign mem[8068] = 5'h11;
  assign mem[8069] = 5'h10;
  assign mem[8070] = 5'h00;
  assign mem[8071] = 5'h01;
  assign mem[8072] = 5'h10;
  assign mem[8073] = 5'h00;
  assign mem[8074] = 5'h02;
  assign mem[8075] = 5'h11;
  assign mem[8076] = 5'h10;
  assign mem[8077] = 5'h00;
  assign mem[8078] = 5'h01;
  assign mem[8079] = 5'h10;
  assign mem[8080] = 5'h00;
  assign mem[8081] = 5'h03;
  assign mem[8082] = 5'h12;
  assign mem[8083] = 5'h11;
  assign mem[8084] = 5'h10;
  assign mem[8085] = 5'h00;
  assign mem[8086] = 5'h01;
  assign mem[8087] = 5'h10;
  assign mem[8088] = 5'h00;
  assign mem[8089] = 5'h02;
  assign mem[8090] = 5'h11;
  assign mem[8091] = 5'h10;
  assign mem[8092] = 5'h00;
  assign mem[8093] = 5'h01;
  assign mem[8094] = 5'h10;
  assign mem[8095] = 5'h00;
  assign mem[8096] = 5'h04;
  assign mem[8097] = 5'h13;
  assign mem[8098] = 5'h12;
  assign mem[8099] = 5'h11;
  assign mem[8100] = 5'h10;
  assign mem[8101] = 5'h00;
  assign mem[8102] = 5'h01;
  assign mem[8103] = 5'h10;
  assign mem[8104] = 5'h00;
  assign mem[8105] = 5'h02;
  assign mem[8106] = 5'h11;
  assign mem[8107] = 5'h10;
  assign mem[8108] = 5'h00;
  assign mem[8109] = 5'h01;
  assign mem[8110] = 5'h10;
  assign mem[8111] = 5'h00;
  assign mem[8112] = 5'h03;
  assign mem[8113] = 5'h12;
  assign mem[8114] = 5'h11;
  assign mem[8115] = 5'h10;
  assign mem[8116] = 5'h00;
  assign mem[8117] = 5'h01;
  assign mem[8118] = 5'h10;
  assign mem[8119] = 5'h00;
  assign mem[8120] = 5'h02;
  assign mem[8121] = 5'h11;
  assign mem[8122] = 5'h10;
  assign mem[8123] = 5'h00;
  assign mem[8124] = 5'h01;
  assign mem[8125] = 5'h10;
  assign mem[8126] = 5'h00;
  assign mem[8127] = 5'h05;
  assign mem[8128] = 5'h14;
  assign mem[8129] = 5'h13;
  assign mem[8130] = 5'h12;
  assign mem[8131] = 5'h11;
  assign mem[8132] = 5'h10;
  assign mem[8133] = 5'h00;
  assign mem[8134] = 5'h01;
  assign mem[8135] = 5'h10;
  assign mem[8136] = 5'h00;
  assign mem[8137] = 5'h02;
  assign mem[8138] = 5'h11;
  assign mem[8139] = 5'h10;
  assign mem[8140] = 5'h00;
  assign mem[8141] = 5'h01;
  assign mem[8142] = 5'h10;
  assign mem[8143] = 5'h00;
  assign mem[8144] = 5'h03;
  assign mem[8145] = 5'h12;
  assign mem[8146] = 5'h11;
  assign mem[8147] = 5'h10;
  assign mem[8148] = 5'h00;
  assign mem[8149] = 5'h01;
  assign mem[8150] = 5'h10;
  assign mem[8151] = 5'h00;
  assign mem[8152] = 5'h02;
  assign mem[8153] = 5'h11;
  assign mem[8154] = 5'h10;
  assign mem[8155] = 5'h00;
  assign mem[8156] = 5'h01;
  assign mem[8157] = 5'h10;
  assign mem[8158] = 5'h00;
  assign mem[8159] = 5'h04;
  assign mem[8160] = 5'h13;
  assign mem[8161] = 5'h12;
  assign mem[8162] = 5'h11;
  assign mem[8163] = 5'h10;
  assign mem[8164] = 5'h00;
  assign mem[8165] = 5'h01;
  assign mem[8166] = 5'h10;
  assign mem[8167] = 5'h00;
  assign mem[8168] = 5'h02;
  assign mem[8169] = 5'h11;
  assign mem[8170] = 5'h10;
  assign mem[8171] = 5'h00;
  assign mem[8172] = 5'h01;
  assign mem[8173] = 5'h10;
  assign mem[8174] = 5'h00;
  assign mem[8175] = 5'h03;
  assign mem[8176] = 5'h12;
  assign mem[8177] = 5'h11;
  assign mem[8178] = 5'h10;
  assign mem[8179] = 5'h00;
  assign mem[8180] = 5'h01;
  assign mem[8181] = 5'h10;
  assign mem[8182] = 5'h00;
  assign mem[8183] = 5'h02;
  assign mem[8184] = 5'h11;
  assign mem[8185] = 5'h10;
  assign mem[8186] = 5'h00;
  assign mem[8187] = 5'h01;
  assign mem[8188] = 5'h10;
  assign mem[8189] = 5'h00;  
  //----
  generate 
  if (RD_TYPE==0)
  begin:U_type0
    reg [$clog2(D)-1:0]addr_d1;

    always @(posedge clk)
    begin
      if((!we) & ce)
        addr_d1 <= addr;
    end

    assign rdata = mem[addr_d1];
  end
  else 
  begin:U_type1

    reg [W-1:0]rdata_int;
    always @(posedge clk)
    begin
      if((!we) & ce)
        rdata_int <= mem[addr];
    end

    assign rdata = rdata_int;
  end
  endgenerate
endmodule
