//////////////////////////////////////////////////////////////////////////////////
// Description:
//////////////////////////////////////////////////////////////////////////////////

module pdec_rom_depth_bd
#(parameter D=16384,
  parameter W=32,
  parameter RD_TYPE=0) //0=delay address by 1T;1=delay rdata
(
  input                 clk,
  input                 ce,   //high active
  input                 we,   //high active
  input  [$clog2(D)-1:0]addr,
  input  [W-1:0]        wdata,
  output [W-1:0]        rdata
);

  wire [W-1:0] mem[0:D-1];
  //----initial
  assign mem[0   ] = 4'h0; 
  assign mem[1   ] = 4'h1;
  assign mem[2   ] = 4'h0;
  assign mem[3   ] = 4'h2;
  assign mem[4   ] = 4'h0;
  assign mem[5   ] = 4'h1;
  assign mem[6   ] = 4'h0;
  assign mem[7   ] = 4'h3;
  assign mem[8   ] = 4'h0;
  assign mem[9   ] = 4'h1;
  assign mem[10  ] = 4'h0;
  assign mem[11  ] = 4'h2;
  assign mem[12  ] = 4'h0;
  assign mem[13  ] = 4'h1;
  assign mem[14  ] = 4'h0;
  assign mem[15  ] = 4'h4;
  assign mem[16  ] = 4'h0;
  assign mem[17  ] = 4'h1;
  assign mem[18  ] = 4'h0;
  assign mem[19  ] = 4'h2;
  assign mem[20  ] = 4'h0;
  assign mem[21  ] = 4'h1;
  assign mem[22  ] = 4'h0;
  assign mem[23  ] = 4'h3;
  assign mem[24  ] = 4'h0;
  assign mem[25  ] = 4'h1;
  assign mem[26  ] = 4'h0;
  assign mem[27  ] = 4'h2;
  assign mem[28  ] = 4'h0;
  assign mem[29  ] = 4'h1;
  assign mem[30  ] = 4'h0;
  assign mem[31  ] = 4'h5;
  assign mem[32  ] = 4'h0;
  assign mem[33  ] = 4'h1;
  assign mem[34  ] = 4'h0;
  assign mem[35  ] = 4'h2;
  assign mem[36  ] = 4'h0;
  assign mem[37  ] = 4'h1;
  assign mem[38  ] = 4'h0;
  assign mem[39  ] = 4'h3;
  assign mem[40  ] = 4'h0;
  assign mem[41  ] = 4'h1;
  assign mem[42  ] = 4'h0;
  assign mem[43  ] = 4'h2;
  assign mem[44  ] = 4'h0;
  assign mem[45  ] = 4'h1;
  assign mem[46  ] = 4'h0;
  assign mem[47  ] = 4'h4;
  assign mem[48  ] = 4'h0;
  assign mem[49  ] = 4'h1;
  assign mem[50  ] = 4'h0;
  assign mem[51  ] = 4'h2;
  assign mem[52  ] = 4'h0;
  assign mem[53  ] = 4'h1;
  assign mem[54  ] = 4'h0;
  assign mem[55  ] = 4'h3;
  assign mem[56  ] = 4'h0;
  assign mem[57  ] = 4'h1;
  assign mem[58  ] = 4'h0;
  assign mem[59  ] = 4'h2;
  assign mem[60  ] = 4'h0;
  assign mem[61  ] = 4'h1;
  assign mem[62  ] = 4'h0;
  assign mem[63  ] = 4'h6;
  assign mem[64  ] = 4'h0;
  assign mem[65  ] = 4'h1;
  assign mem[66  ] = 4'h0;
  assign mem[67  ] = 4'h2;
  assign mem[68  ] = 4'h0;
  assign mem[69  ] = 4'h1;
  assign mem[70  ] = 4'h0;
  assign mem[71  ] = 4'h3;
  assign mem[72  ] = 4'h0;
  assign mem[73  ] = 4'h1;
  assign mem[74  ] = 4'h0;
  assign mem[75  ] = 4'h2;
  assign mem[76  ] = 4'h0;
  assign mem[77  ] = 4'h1;
  assign mem[78  ] = 4'h0;
  assign mem[79  ] = 4'h4;
  assign mem[80  ] = 4'h0;
  assign mem[81  ] = 4'h1;
  assign mem[82  ] = 4'h0;
  assign mem[83  ] = 4'h2;
  assign mem[84  ] = 4'h0;
  assign mem[85  ] = 4'h1;
  assign mem[86  ] = 4'h0;
  assign mem[87  ] = 4'h3;
  assign mem[88  ] = 4'h0;
  assign mem[89  ] = 4'h1;
  assign mem[90  ] = 4'h0;
  assign mem[91  ] = 4'h2;
  assign mem[92  ] = 4'h0;
  assign mem[93  ] = 4'h1;
  assign mem[94  ] = 4'h0;
  assign mem[95  ] = 4'h5;
  assign mem[96  ] = 4'h0;
  assign mem[97  ] = 4'h1;
  assign mem[98  ] = 4'h0;
  assign mem[99  ] = 4'h2;
  assign mem[100 ] = 4'h0;
  assign mem[101 ] = 4'h1;
  assign mem[102 ] = 4'h0;
  assign mem[103 ] = 4'h3;
  assign mem[104 ] = 4'h0;
  assign mem[105 ] = 4'h1;
  assign mem[106 ] = 4'h0;
  assign mem[107 ] = 4'h2;
  assign mem[108 ] = 4'h0;
  assign mem[109 ] = 4'h1;
  assign mem[110 ] = 4'h0;
  assign mem[111 ] = 4'h4;
  assign mem[112 ] = 4'h0;
  assign mem[113 ] = 4'h1;
  assign mem[114 ] = 4'h0;
  assign mem[115 ] = 4'h2;
  assign mem[116 ] = 4'h0;
  assign mem[117 ] = 4'h1;
  assign mem[118 ] = 4'h0;
  assign mem[119 ] = 4'h3;
  assign mem[120 ] = 4'h0;
  assign mem[121 ] = 4'h1;
  assign mem[122 ] = 4'h0;
  assign mem[123 ] = 4'h2;
  assign mem[124 ] = 4'h0;
  assign mem[125 ] = 4'h1;
  assign mem[126 ] = 4'h0;
  assign mem[127 ] = 4'h7;
  assign mem[128 ] = 4'h0;
  assign mem[129 ] = 4'h1;
  assign mem[130 ] = 4'h0;
  assign mem[131 ] = 4'h2;
  assign mem[132 ] = 4'h0;
  assign mem[133 ] = 4'h1;
  assign mem[134 ] = 4'h0;
  assign mem[135 ] = 4'h3;
  assign mem[136 ] = 4'h0;
  assign mem[137 ] = 4'h1;
  assign mem[138 ] = 4'h0;
  assign mem[139 ] = 4'h2;
  assign mem[140 ] = 4'h0;
  assign mem[141 ] = 4'h1;
  assign mem[142 ] = 4'h0;
  assign mem[143 ] = 4'h4;
  assign mem[144 ] = 4'h0;
  assign mem[145 ] = 4'h1;
  assign mem[146 ] = 4'h0;
  assign mem[147 ] = 4'h2;
  assign mem[148 ] = 4'h0;
  assign mem[149 ] = 4'h1;
  assign mem[150 ] = 4'h0;
  assign mem[151 ] = 4'h3;
  assign mem[152 ] = 4'h0;
  assign mem[153 ] = 4'h1;
  assign mem[154 ] = 4'h0;
  assign mem[155 ] = 4'h2;
  assign mem[156 ] = 4'h0;
  assign mem[157 ] = 4'h1;
  assign mem[158 ] = 4'h0;
  assign mem[159 ] = 4'h5;
  assign mem[160 ] = 4'h0;
  assign mem[161 ] = 4'h1;
  assign mem[162 ] = 4'h0;
  assign mem[163 ] = 4'h2;
  assign mem[164 ] = 4'h0;
  assign mem[165 ] = 4'h1;
  assign mem[166 ] = 4'h0;
  assign mem[167 ] = 4'h3;
  assign mem[168 ] = 4'h0;
  assign mem[169 ] = 4'h1;
  assign mem[170 ] = 4'h0;
  assign mem[171 ] = 4'h2;
  assign mem[172 ] = 4'h0;
  assign mem[173 ] = 4'h1;
  assign mem[174 ] = 4'h0;
  assign mem[175 ] = 4'h4;
  assign mem[176 ] = 4'h0;
  assign mem[177 ] = 4'h1;
  assign mem[178 ] = 4'h0;
  assign mem[179 ] = 4'h2;
  assign mem[180 ] = 4'h0;
  assign mem[181 ] = 4'h1;
  assign mem[182 ] = 4'h0;
  assign mem[183 ] = 4'h3;
  assign mem[184 ] = 4'h0;
  assign mem[185 ] = 4'h1;
  assign mem[186 ] = 4'h0;
  assign mem[187 ] = 4'h2;
  assign mem[188 ] = 4'h0;
  assign mem[189 ] = 4'h1;
  assign mem[190 ] = 4'h0;
  assign mem[191 ] = 4'h6;
  assign mem[192 ] = 4'h0;
  assign mem[193 ] = 4'h1;
  assign mem[194 ] = 4'h0;
  assign mem[195 ] = 4'h2;
  assign mem[196 ] = 4'h0;
  assign mem[197 ] = 4'h1;
  assign mem[198 ] = 4'h0;
  assign mem[199 ] = 4'h3;
  assign mem[200 ] = 4'h0;
  assign mem[201 ] = 4'h1;
  assign mem[202 ] = 4'h0;
  assign mem[203 ] = 4'h2;
  assign mem[204 ] = 4'h0;
  assign mem[205 ] = 4'h1;
  assign mem[206 ] = 4'h0;
  assign mem[207 ] = 4'h4;
  assign mem[208 ] = 4'h0;
  assign mem[209 ] = 4'h1;
  assign mem[210 ] = 4'h0;
  assign mem[211 ] = 4'h2;
  assign mem[212 ] = 4'h0;
  assign mem[213 ] = 4'h1;
  assign mem[214 ] = 4'h0;
  assign mem[215 ] = 4'h3;
  assign mem[216 ] = 4'h0;
  assign mem[217 ] = 4'h1;
  assign mem[218 ] = 4'h0;
  assign mem[219 ] = 4'h2;
  assign mem[220 ] = 4'h0;
  assign mem[221 ] = 4'h1;
  assign mem[222 ] = 4'h0;
  assign mem[223 ] = 4'h5;
  assign mem[224 ] = 4'h0;
  assign mem[225 ] = 4'h1;
  assign mem[226 ] = 4'h0;
  assign mem[227 ] = 4'h2;
  assign mem[228 ] = 4'h0;
  assign mem[229 ] = 4'h1;
  assign mem[230 ] = 4'h0;
  assign mem[231 ] = 4'h3;
  assign mem[232 ] = 4'h0;
  assign mem[233 ] = 4'h1;
  assign mem[234 ] = 4'h0;
  assign mem[235 ] = 4'h2;
  assign mem[236 ] = 4'h0;
  assign mem[237 ] = 4'h1;
  assign mem[238 ] = 4'h0;
  assign mem[239 ] = 4'h4;
  assign mem[240 ] = 4'h0;
  assign mem[241 ] = 4'h1;
  assign mem[242 ] = 4'h0;
  assign mem[243 ] = 4'h2;
  assign mem[244 ] = 4'h0;
  assign mem[245 ] = 4'h1;
  assign mem[246 ] = 4'h0;
  assign mem[247 ] = 4'h3;
  assign mem[248 ] = 4'h0;
  assign mem[249 ] = 4'h1;
  assign mem[250 ] = 4'h0;
  assign mem[251 ] = 4'h2;
  assign mem[252 ] = 4'h0;
  assign mem[253 ] = 4'h1;
  assign mem[254 ] = 4'h0;
  assign mem[255 ] = 4'h8;
  assign mem[256 ] = 4'h0;
  assign mem[257 ] = 4'h1;
  assign mem[258 ] = 4'h0;
  assign mem[259 ] = 4'h2;
  assign mem[260 ] = 4'h0;
  assign mem[261 ] = 4'h1;
  assign mem[262 ] = 4'h0;
  assign mem[263 ] = 4'h3;
  assign mem[264 ] = 4'h0;
  assign mem[265 ] = 4'h1;
  assign mem[266 ] = 4'h0;
  assign mem[267 ] = 4'h2;
  assign mem[268 ] = 4'h0;
  assign mem[269 ] = 4'h1;
  assign mem[270 ] = 4'h0;
  assign mem[271 ] = 4'h4;
  assign mem[272 ] = 4'h0;
  assign mem[273 ] = 4'h1;
  assign mem[274 ] = 4'h0;
  assign mem[275 ] = 4'h2;
  assign mem[276 ] = 4'h0;
  assign mem[277 ] = 4'h1;
  assign mem[278 ] = 4'h0;
  assign mem[279 ] = 4'h3;
  assign mem[280 ] = 4'h0;
  assign mem[281 ] = 4'h1;
  assign mem[282 ] = 4'h0;
  assign mem[283 ] = 4'h2;
  assign mem[284 ] = 4'h0;
  assign mem[285 ] = 4'h1;
  assign mem[286 ] = 4'h0;
  assign mem[287 ] = 4'h5;
  assign mem[288 ] = 4'h0;
  assign mem[289 ] = 4'h1;
  assign mem[290 ] = 4'h0;
  assign mem[291 ] = 4'h2;
  assign mem[292 ] = 4'h0;
  assign mem[293 ] = 4'h1;
  assign mem[294 ] = 4'h0;
  assign mem[295 ] = 4'h3;
  assign mem[296 ] = 4'h0;
  assign mem[297 ] = 4'h1;
  assign mem[298 ] = 4'h0;
  assign mem[299 ] = 4'h2;
  assign mem[300 ] = 4'h0;
  assign mem[301 ] = 4'h1;
  assign mem[302 ] = 4'h0;
  assign mem[303 ] = 4'h4;
  assign mem[304 ] = 4'h0;
  assign mem[305 ] = 4'h1;
  assign mem[306 ] = 4'h0;
  assign mem[307 ] = 4'h2;
  assign mem[308 ] = 4'h0;
  assign mem[309 ] = 4'h1;
  assign mem[310 ] = 4'h0;
  assign mem[311 ] = 4'h3;
  assign mem[312 ] = 4'h0;
  assign mem[313 ] = 4'h1;
  assign mem[314 ] = 4'h0;
  assign mem[315 ] = 4'h2;
  assign mem[316 ] = 4'h0;
  assign mem[317 ] = 4'h1;
  assign mem[318 ] = 4'h0;
  assign mem[319 ] = 4'h6;
  assign mem[320 ] = 4'h0;
  assign mem[321 ] = 4'h1;
  assign mem[322 ] = 4'h0;
  assign mem[323 ] = 4'h2;
  assign mem[324 ] = 4'h0;
  assign mem[325 ] = 4'h1;
  assign mem[326 ] = 4'h0;
  assign mem[327 ] = 4'h3;
  assign mem[328 ] = 4'h0;
  assign mem[329 ] = 4'h1;
  assign mem[330 ] = 4'h0;
  assign mem[331 ] = 4'h2;
  assign mem[332 ] = 4'h0;
  assign mem[333 ] = 4'h1;
  assign mem[334 ] = 4'h0;
  assign mem[335 ] = 4'h4;
  assign mem[336 ] = 4'h0;
  assign mem[337 ] = 4'h1;
  assign mem[338 ] = 4'h0;
  assign mem[339 ] = 4'h2;
  assign mem[340 ] = 4'h0;
  assign mem[341 ] = 4'h1;
  assign mem[342 ] = 4'h0;
  assign mem[343 ] = 4'h3;
  assign mem[344 ] = 4'h0;
  assign mem[345 ] = 4'h1;
  assign mem[346 ] = 4'h0;
  assign mem[347 ] = 4'h2;
  assign mem[348 ] = 4'h0;
  assign mem[349 ] = 4'h1;
  assign mem[350 ] = 4'h0;
  assign mem[351 ] = 4'h5;
  assign mem[352 ] = 4'h0;
  assign mem[353 ] = 4'h1;
  assign mem[354 ] = 4'h0;
  assign mem[355 ] = 4'h2;
  assign mem[356 ] = 4'h0;
  assign mem[357 ] = 4'h1;
  assign mem[358 ] = 4'h0;
  assign mem[359 ] = 4'h3;
  assign mem[360 ] = 4'h0;
  assign mem[361 ] = 4'h1;
  assign mem[362 ] = 4'h0;
  assign mem[363 ] = 4'h2;
  assign mem[364 ] = 4'h0;
  assign mem[365 ] = 4'h1;
  assign mem[366 ] = 4'h0;
  assign mem[367 ] = 4'h4;
  assign mem[368 ] = 4'h0;
  assign mem[369 ] = 4'h1;
  assign mem[370 ] = 4'h0;
  assign mem[371 ] = 4'h2;
  assign mem[372 ] = 4'h0;
  assign mem[373 ] = 4'h1;
  assign mem[374 ] = 4'h0;
  assign mem[375 ] = 4'h3;
  assign mem[376 ] = 4'h0;
  assign mem[377 ] = 4'h1;
  assign mem[378 ] = 4'h0;
  assign mem[379 ] = 4'h2;
  assign mem[380 ] = 4'h0;
  assign mem[381 ] = 4'h1;
  assign mem[382 ] = 4'h0;
  assign mem[383 ] = 4'h7;
  assign mem[384 ] = 4'h0;
  assign mem[385 ] = 4'h1;
  assign mem[386 ] = 4'h0;
  assign mem[387 ] = 4'h2;
  assign mem[388 ] = 4'h0;
  assign mem[389 ] = 4'h1;
  assign mem[390 ] = 4'h0;
  assign mem[391 ] = 4'h3;
  assign mem[392 ] = 4'h0;
  assign mem[393 ] = 4'h1;
  assign mem[394 ] = 4'h0;
  assign mem[395 ] = 4'h2;
  assign mem[396 ] = 4'h0;
  assign mem[397 ] = 4'h1;
  assign mem[398 ] = 4'h0;
  assign mem[399 ] = 4'h4;
  assign mem[400 ] = 4'h0;
  assign mem[401 ] = 4'h1;
  assign mem[402 ] = 4'h0;
  assign mem[403 ] = 4'h2;
  assign mem[404 ] = 4'h0;
  assign mem[405 ] = 4'h1;
  assign mem[406 ] = 4'h0;
  assign mem[407 ] = 4'h3;
  assign mem[408 ] = 4'h0;
  assign mem[409 ] = 4'h1;
  assign mem[410 ] = 4'h0;
  assign mem[411 ] = 4'h2;
  assign mem[412 ] = 4'h0;
  assign mem[413 ] = 4'h1;
  assign mem[414 ] = 4'h0;
  assign mem[415 ] = 4'h5;
  assign mem[416 ] = 4'h0;
  assign mem[417 ] = 4'h1;
  assign mem[418 ] = 4'h0;
  assign mem[419 ] = 4'h2;
  assign mem[420 ] = 4'h0;
  assign mem[421 ] = 4'h1;
  assign mem[422 ] = 4'h0;
  assign mem[423 ] = 4'h3;
  assign mem[424 ] = 4'h0;
  assign mem[425 ] = 4'h1;
  assign mem[426 ] = 4'h0;
  assign mem[427 ] = 4'h2;
  assign mem[428 ] = 4'h0;
  assign mem[429 ] = 4'h1;
  assign mem[430 ] = 4'h0;
  assign mem[431 ] = 4'h4;
  assign mem[432 ] = 4'h0;
  assign mem[433 ] = 4'h1;
  assign mem[434 ] = 4'h0;
  assign mem[435 ] = 4'h2;
  assign mem[436 ] = 4'h0;
  assign mem[437 ] = 4'h1;
  assign mem[438 ] = 4'h0;
  assign mem[439 ] = 4'h3;
  assign mem[440 ] = 4'h0;
  assign mem[441 ] = 4'h1;
  assign mem[442 ] = 4'h0;
  assign mem[443 ] = 4'h2;
  assign mem[444 ] = 4'h0;
  assign mem[445 ] = 4'h1;
  assign mem[446 ] = 4'h0;
  assign mem[447 ] = 4'h6;
  assign mem[448 ] = 4'h0;
  assign mem[449 ] = 4'h1;
  assign mem[450 ] = 4'h0;
  assign mem[451 ] = 4'h2;
  assign mem[452 ] = 4'h0;
  assign mem[453 ] = 4'h1;
  assign mem[454 ] = 4'h0;
  assign mem[455 ] = 4'h3;
  assign mem[456 ] = 4'h0;
  assign mem[457 ] = 4'h1;
  assign mem[458 ] = 4'h0;
  assign mem[459 ] = 4'h2;
  assign mem[460 ] = 4'h0;
  assign mem[461 ] = 4'h1;
  assign mem[462 ] = 4'h0;
  assign mem[463 ] = 4'h4;
  assign mem[464 ] = 4'h0;
  assign mem[465 ] = 4'h1;
  assign mem[466 ] = 4'h0;
  assign mem[467 ] = 4'h2;
  assign mem[468 ] = 4'h0;
  assign mem[469 ] = 4'h1;
  assign mem[470 ] = 4'h0;
  assign mem[471 ] = 4'h3;
  assign mem[472 ] = 4'h0;
  assign mem[473 ] = 4'h1;
  assign mem[474 ] = 4'h0;
  assign mem[475 ] = 4'h2;
  assign mem[476 ] = 4'h0;
  assign mem[477 ] = 4'h1;
  assign mem[478 ] = 4'h0;
  assign mem[479 ] = 4'h5;
  assign mem[480 ] = 4'h0;
  assign mem[481 ] = 4'h1;
  assign mem[482 ] = 4'h0;
  assign mem[483 ] = 4'h2;
  assign mem[484 ] = 4'h0;
  assign mem[485 ] = 4'h1;
  assign mem[486 ] = 4'h0;
  assign mem[487 ] = 4'h3;
  assign mem[488 ] = 4'h0;
  assign mem[489 ] = 4'h1;
  assign mem[490 ] = 4'h0;
  assign mem[491 ] = 4'h2;
  assign mem[492 ] = 4'h0;
  assign mem[493 ] = 4'h1;
  assign mem[494 ] = 4'h0;
  assign mem[495 ] = 4'h4;
  assign mem[496 ] = 4'h0;
  assign mem[497 ] = 4'h1;
  assign mem[498 ] = 4'h0;
  assign mem[499 ] = 4'h2;
  assign mem[500 ] = 4'h0;
  assign mem[501 ] = 4'h1;
  assign mem[502 ] = 4'h0;
  assign mem[503 ] = 4'h3;
  assign mem[504 ] = 4'h0;
  assign mem[505 ] = 4'h1;
  assign mem[506 ] = 4'h0;
  assign mem[507 ] = 4'h2;
  assign mem[508 ] = 4'h0;
  assign mem[509 ] = 4'h1;
  assign mem[510 ] = 4'h0;
  assign mem[511 ] = 4'h9;
  assign mem[512 ] = 4'h0;
  assign mem[513 ] = 4'h1;
  assign mem[514 ] = 4'h0;
  assign mem[515 ] = 4'h2;
  assign mem[516 ] = 4'h0;
  assign mem[517 ] = 4'h1;
  assign mem[518 ] = 4'h0;
  assign mem[519 ] = 4'h3;
  assign mem[520 ] = 4'h0;
  assign mem[521 ] = 4'h1;
  assign mem[522 ] = 4'h0;
  assign mem[523 ] = 4'h2;
  assign mem[524 ] = 4'h0;
  assign mem[525 ] = 4'h1;
  assign mem[526 ] = 4'h0;
  assign mem[527 ] = 4'h4;
  assign mem[528 ] = 4'h0;
  assign mem[529 ] = 4'h1;
  assign mem[530 ] = 4'h0;
  assign mem[531 ] = 4'h2;
  assign mem[532 ] = 4'h0;
  assign mem[533 ] = 4'h1;
  assign mem[534 ] = 4'h0;
  assign mem[535 ] = 4'h3;
  assign mem[536 ] = 4'h0;
  assign mem[537 ] = 4'h1;
  assign mem[538 ] = 4'h0;
  assign mem[539 ] = 4'h2;
  assign mem[540 ] = 4'h0;
  assign mem[541 ] = 4'h1;
  assign mem[542 ] = 4'h0;
  assign mem[543 ] = 4'h5;
  assign mem[544 ] = 4'h0;
  assign mem[545 ] = 4'h1;
  assign mem[546 ] = 4'h0;
  assign mem[547 ] = 4'h2;
  assign mem[548 ] = 4'h0;
  assign mem[549 ] = 4'h1;
  assign mem[550 ] = 4'h0;
  assign mem[551 ] = 4'h3;
  assign mem[552 ] = 4'h0;
  assign mem[553 ] = 4'h1;
  assign mem[554 ] = 4'h0;
  assign mem[555 ] = 4'h2;
  assign mem[556 ] = 4'h0;
  assign mem[557 ] = 4'h1;
  assign mem[558 ] = 4'h0;
  assign mem[559 ] = 4'h4;
  assign mem[560 ] = 4'h0;
  assign mem[561 ] = 4'h1;
  assign mem[562 ] = 4'h0;
  assign mem[563 ] = 4'h2;
  assign mem[564 ] = 4'h0;
  assign mem[565 ] = 4'h1;
  assign mem[566 ] = 4'h0;
  assign mem[567 ] = 4'h3;
  assign mem[568 ] = 4'h0;
  assign mem[569 ] = 4'h1;
  assign mem[570 ] = 4'h0;
  assign mem[571 ] = 4'h2;
  assign mem[572 ] = 4'h0;
  assign mem[573 ] = 4'h1;
  assign mem[574 ] = 4'h0;
  assign mem[575 ] = 4'h6;
  assign mem[576 ] = 4'h0;
  assign mem[577 ] = 4'h1;
  assign mem[578 ] = 4'h0;
  assign mem[579 ] = 4'h2;
  assign mem[580 ] = 4'h0;
  assign mem[581 ] = 4'h1;
  assign mem[582 ] = 4'h0;
  assign mem[583 ] = 4'h3;
  assign mem[584 ] = 4'h0;
  assign mem[585 ] = 4'h1;
  assign mem[586 ] = 4'h0;
  assign mem[587 ] = 4'h2;
  assign mem[588 ] = 4'h0;
  assign mem[589 ] = 4'h1;
  assign mem[590 ] = 4'h0;
  assign mem[591 ] = 4'h4;
  assign mem[592 ] = 4'h0;
  assign mem[593 ] = 4'h1;
  assign mem[594 ] = 4'h0;
  assign mem[595 ] = 4'h2;
  assign mem[596 ] = 4'h0;
  assign mem[597 ] = 4'h1;
  assign mem[598 ] = 4'h0;
  assign mem[599 ] = 4'h3;
  assign mem[600 ] = 4'h0;
  assign mem[601 ] = 4'h1;
  assign mem[602 ] = 4'h0;
  assign mem[603 ] = 4'h2;
  assign mem[604 ] = 4'h0;
  assign mem[605 ] = 4'h1;
  assign mem[606 ] = 4'h0;
  assign mem[607 ] = 4'h5;
  assign mem[608 ] = 4'h0;
  assign mem[609 ] = 4'h1;
  assign mem[610 ] = 4'h0;
  assign mem[611 ] = 4'h2;
  assign mem[612 ] = 4'h0;
  assign mem[613 ] = 4'h1;
  assign mem[614 ] = 4'h0;
  assign mem[615 ] = 4'h3;
  assign mem[616 ] = 4'h0;
  assign mem[617 ] = 4'h1;
  assign mem[618 ] = 4'h0;
  assign mem[619 ] = 4'h2;
  assign mem[620 ] = 4'h0;
  assign mem[621 ] = 4'h1;
  assign mem[622 ] = 4'h0;
  assign mem[623 ] = 4'h4;
  assign mem[624 ] = 4'h0;
  assign mem[625 ] = 4'h1;
  assign mem[626 ] = 4'h0;
  assign mem[627 ] = 4'h2;
  assign mem[628 ] = 4'h0;
  assign mem[629 ] = 4'h1;
  assign mem[630 ] = 4'h0;
  assign mem[631 ] = 4'h3;
  assign mem[632 ] = 4'h0;
  assign mem[633 ] = 4'h1;
  assign mem[634 ] = 4'h0;
  assign mem[635 ] = 4'h2;
  assign mem[636 ] = 4'h0;
  assign mem[637 ] = 4'h1;
  assign mem[638 ] = 4'h0;
  assign mem[639 ] = 4'h7;
  assign mem[640 ] = 4'h0;
  assign mem[641 ] = 4'h1;
  assign mem[642 ] = 4'h0;
  assign mem[643 ] = 4'h2;
  assign mem[644 ] = 4'h0;
  assign mem[645 ] = 4'h1;
  assign mem[646 ] = 4'h0;
  assign mem[647 ] = 4'h3;
  assign mem[648 ] = 4'h0;
  assign mem[649 ] = 4'h1;
  assign mem[650 ] = 4'h0;
  assign mem[651 ] = 4'h2;
  assign mem[652 ] = 4'h0;
  assign mem[653 ] = 4'h1;
  assign mem[654 ] = 4'h0;
  assign mem[655 ] = 4'h4;
  assign mem[656 ] = 4'h0;
  assign mem[657 ] = 4'h1;
  assign mem[658 ] = 4'h0;
  assign mem[659 ] = 4'h2;
  assign mem[660 ] = 4'h0;
  assign mem[661 ] = 4'h1;
  assign mem[662 ] = 4'h0;
  assign mem[663 ] = 4'h3;
  assign mem[664 ] = 4'h0;
  assign mem[665 ] = 4'h1;
  assign mem[666 ] = 4'h0;
  assign mem[667 ] = 4'h2;
  assign mem[668 ] = 4'h0;
  assign mem[669 ] = 4'h1;
  assign mem[670 ] = 4'h0;
  assign mem[671 ] = 4'h5;
  assign mem[672 ] = 4'h0;
  assign mem[673 ] = 4'h1;
  assign mem[674 ] = 4'h0;
  assign mem[675 ] = 4'h2;
  assign mem[676 ] = 4'h0;
  assign mem[677 ] = 4'h1;
  assign mem[678 ] = 4'h0;
  assign mem[679 ] = 4'h3;
  assign mem[680 ] = 4'h0;
  assign mem[681 ] = 4'h1;
  assign mem[682 ] = 4'h0;
  assign mem[683 ] = 4'h2;
  assign mem[684 ] = 4'h0;
  assign mem[685 ] = 4'h1;
  assign mem[686 ] = 4'h0;
  assign mem[687 ] = 4'h4;
  assign mem[688 ] = 4'h0;
  assign mem[689 ] = 4'h1;
  assign mem[690 ] = 4'h0;
  assign mem[691 ] = 4'h2;
  assign mem[692 ] = 4'h0;
  assign mem[693 ] = 4'h1;
  assign mem[694 ] = 4'h0;
  assign mem[695 ] = 4'h3;
  assign mem[696 ] = 4'h0;
  assign mem[697 ] = 4'h1;
  assign mem[698 ] = 4'h0;
  assign mem[699 ] = 4'h2;
  assign mem[700 ] = 4'h0;
  assign mem[701 ] = 4'h1;
  assign mem[702 ] = 4'h0;
  assign mem[703 ] = 4'h6;
  assign mem[704 ] = 4'h0;
  assign mem[705 ] = 4'h1;
  assign mem[706 ] = 4'h0;
  assign mem[707 ] = 4'h2;
  assign mem[708 ] = 4'h0;
  assign mem[709 ] = 4'h1;
  assign mem[710 ] = 4'h0;
  assign mem[711 ] = 4'h3;
  assign mem[712 ] = 4'h0;
  assign mem[713 ] = 4'h1;
  assign mem[714 ] = 4'h0;
  assign mem[715 ] = 4'h2;
  assign mem[716 ] = 4'h0;
  assign mem[717 ] = 4'h1;
  assign mem[718 ] = 4'h0;
  assign mem[719 ] = 4'h4;
  assign mem[720 ] = 4'h0;
  assign mem[721 ] = 4'h1;
  assign mem[722 ] = 4'h0;
  assign mem[723 ] = 4'h2;
  assign mem[724 ] = 4'h0;
  assign mem[725 ] = 4'h1;
  assign mem[726 ] = 4'h0;
  assign mem[727 ] = 4'h3;
  assign mem[728 ] = 4'h0;
  assign mem[729 ] = 4'h1;
  assign mem[730 ] = 4'h0;
  assign mem[731 ] = 4'h2;
  assign mem[732 ] = 4'h0;
  assign mem[733 ] = 4'h1;
  assign mem[734 ] = 4'h0;
  assign mem[735 ] = 4'h5;
  assign mem[736 ] = 4'h0;
  assign mem[737 ] = 4'h1;
  assign mem[738 ] = 4'h0;
  assign mem[739 ] = 4'h2;
  assign mem[740 ] = 4'h0;
  assign mem[741 ] = 4'h1;
  assign mem[742 ] = 4'h0;
  assign mem[743 ] = 4'h3;
  assign mem[744 ] = 4'h0;
  assign mem[745 ] = 4'h1;
  assign mem[746 ] = 4'h0;
  assign mem[747 ] = 4'h2;
  assign mem[748 ] = 4'h0;
  assign mem[749 ] = 4'h1;
  assign mem[750 ] = 4'h0;
  assign mem[751 ] = 4'h4;
  assign mem[752 ] = 4'h0;
  assign mem[753 ] = 4'h1;
  assign mem[754 ] = 4'h0;
  assign mem[755 ] = 4'h2;
  assign mem[756 ] = 4'h0;
  assign mem[757 ] = 4'h1;
  assign mem[758 ] = 4'h0;
  assign mem[759 ] = 4'h3;
  assign mem[760 ] = 4'h0;
  assign mem[761 ] = 4'h1;
  assign mem[762 ] = 4'h0;
  assign mem[763 ] = 4'h2;
  assign mem[764 ] = 4'h0;
  assign mem[765 ] = 4'h1;
  assign mem[766 ] = 4'h0;
  assign mem[767 ] = 4'h8;
  assign mem[768 ] = 4'h0;
  assign mem[769 ] = 4'h1;
  assign mem[770 ] = 4'h0;
  assign mem[771 ] = 4'h2;
  assign mem[772 ] = 4'h0;
  assign mem[773 ] = 4'h1;
  assign mem[774 ] = 4'h0;
  assign mem[775 ] = 4'h3;
  assign mem[776 ] = 4'h0;
  assign mem[777 ] = 4'h1;
  assign mem[778 ] = 4'h0;
  assign mem[779 ] = 4'h2;
  assign mem[780 ] = 4'h0;
  assign mem[781 ] = 4'h1;
  assign mem[782 ] = 4'h0;
  assign mem[783 ] = 4'h4;
  assign mem[784 ] = 4'h0;
  assign mem[785 ] = 4'h1;
  assign mem[786 ] = 4'h0;
  assign mem[787 ] = 4'h2;
  assign mem[788 ] = 4'h0;
  assign mem[789 ] = 4'h1;
  assign mem[790 ] = 4'h0;
  assign mem[791 ] = 4'h3;
  assign mem[792 ] = 4'h0;
  assign mem[793 ] = 4'h1;
  assign mem[794 ] = 4'h0;
  assign mem[795 ] = 4'h2;
  assign mem[796 ] = 4'h0;
  assign mem[797 ] = 4'h1;
  assign mem[798 ] = 4'h0;
  assign mem[799 ] = 4'h5;
  assign mem[800 ] = 4'h0;
  assign mem[801 ] = 4'h1;
  assign mem[802 ] = 4'h0;
  assign mem[803 ] = 4'h2;
  assign mem[804 ] = 4'h0;
  assign mem[805 ] = 4'h1;
  assign mem[806 ] = 4'h0;
  assign mem[807 ] = 4'h3;
  assign mem[808 ] = 4'h0;
  assign mem[809 ] = 4'h1;
  assign mem[810 ] = 4'h0;
  assign mem[811 ] = 4'h2;
  assign mem[812 ] = 4'h0;
  assign mem[813 ] = 4'h1;
  assign mem[814 ] = 4'h0;
  assign mem[815 ] = 4'h4;
  assign mem[816 ] = 4'h0;
  assign mem[817 ] = 4'h1;
  assign mem[818 ] = 4'h0;
  assign mem[819 ] = 4'h2;
  assign mem[820 ] = 4'h0;
  assign mem[821 ] = 4'h1;
  assign mem[822 ] = 4'h0;
  assign mem[823 ] = 4'h3;
  assign mem[824 ] = 4'h0;
  assign mem[825 ] = 4'h1;
  assign mem[826 ] = 4'h0;
  assign mem[827 ] = 4'h2;
  assign mem[828 ] = 4'h0;
  assign mem[829 ] = 4'h1;
  assign mem[830 ] = 4'h0;
  assign mem[831 ] = 4'h6;
  assign mem[832 ] = 4'h0;
  assign mem[833 ] = 4'h1;
  assign mem[834 ] = 4'h0;
  assign mem[835 ] = 4'h2;
  assign mem[836 ] = 4'h0;
  assign mem[837 ] = 4'h1;
  assign mem[838 ] = 4'h0;
  assign mem[839 ] = 4'h3;
  assign mem[840 ] = 4'h0;
  assign mem[841 ] = 4'h1;
  assign mem[842 ] = 4'h0;
  assign mem[843 ] = 4'h2;
  assign mem[844 ] = 4'h0;
  assign mem[845 ] = 4'h1;
  assign mem[846 ] = 4'h0;
  assign mem[847 ] = 4'h4;
  assign mem[848 ] = 4'h0;
  assign mem[849 ] = 4'h1;
  assign mem[850 ] = 4'h0;
  assign mem[851 ] = 4'h2;
  assign mem[852 ] = 4'h0;
  assign mem[853 ] = 4'h1;
  assign mem[854 ] = 4'h0;
  assign mem[855 ] = 4'h3;
  assign mem[856 ] = 4'h0;
  assign mem[857 ] = 4'h1;
  assign mem[858 ] = 4'h0;
  assign mem[859 ] = 4'h2;
  assign mem[860 ] = 4'h0;
  assign mem[861 ] = 4'h1;
  assign mem[862 ] = 4'h0;
  assign mem[863 ] = 4'h5;
  assign mem[864 ] = 4'h0;
  assign mem[865 ] = 4'h1;
  assign mem[866 ] = 4'h0;
  assign mem[867 ] = 4'h2;
  assign mem[868 ] = 4'h0;
  assign mem[869 ] = 4'h1;
  assign mem[870 ] = 4'h0;
  assign mem[871 ] = 4'h3;
  assign mem[872 ] = 4'h0;
  assign mem[873 ] = 4'h1;
  assign mem[874 ] = 4'h0;
  assign mem[875 ] = 4'h2;
  assign mem[876 ] = 4'h0;
  assign mem[877 ] = 4'h1;
  assign mem[878 ] = 4'h0;
  assign mem[879 ] = 4'h4;
  assign mem[880 ] = 4'h0;
  assign mem[881 ] = 4'h1;
  assign mem[882 ] = 4'h0;
  assign mem[883 ] = 4'h2;
  assign mem[884 ] = 4'h0;
  assign mem[885 ] = 4'h1;
  assign mem[886 ] = 4'h0;
  assign mem[887 ] = 4'h3;
  assign mem[888 ] = 4'h0;
  assign mem[889 ] = 4'h1;
  assign mem[890 ] = 4'h0;
  assign mem[891 ] = 4'h2;
  assign mem[892 ] = 4'h0;
  assign mem[893 ] = 4'h1;
  assign mem[894 ] = 4'h0;
  assign mem[895 ] = 4'h7;
  assign mem[896 ] = 4'h0;
  assign mem[897 ] = 4'h1;
  assign mem[898 ] = 4'h0;
  assign mem[899 ] = 4'h2;
  assign mem[900 ] = 4'h0;
  assign mem[901 ] = 4'h1;
  assign mem[902 ] = 4'h0;
  assign mem[903 ] = 4'h3;
  assign mem[904 ] = 4'h0;
  assign mem[905 ] = 4'h1;
  assign mem[906 ] = 4'h0;
  assign mem[907 ] = 4'h2;
  assign mem[908 ] = 4'h0;
  assign mem[909 ] = 4'h1;
  assign mem[910 ] = 4'h0;
  assign mem[911 ] = 4'h4;
  assign mem[912 ] = 4'h0;
  assign mem[913 ] = 4'h1;
  assign mem[914 ] = 4'h0;
  assign mem[915 ] = 4'h2;
  assign mem[916 ] = 4'h0;
  assign mem[917 ] = 4'h1;
  assign mem[918 ] = 4'h0;
  assign mem[919 ] = 4'h3;
  assign mem[920 ] = 4'h0;
  assign mem[921 ] = 4'h1;
  assign mem[922 ] = 4'h0;
  assign mem[923 ] = 4'h2;
  assign mem[924 ] = 4'h0;
  assign mem[925 ] = 4'h1;
  assign mem[926 ] = 4'h0;
  assign mem[927 ] = 4'h5;
  assign mem[928 ] = 4'h0;
  assign mem[929 ] = 4'h1;
  assign mem[930 ] = 4'h0;
  assign mem[931 ] = 4'h2;
  assign mem[932 ] = 4'h0;
  assign mem[933 ] = 4'h1;
  assign mem[934 ] = 4'h0;
  assign mem[935 ] = 4'h3;
  assign mem[936 ] = 4'h0;
  assign mem[937 ] = 4'h1;
  assign mem[938 ] = 4'h0;
  assign mem[939 ] = 4'h2;
  assign mem[940 ] = 4'h0;
  assign mem[941 ] = 4'h1;
  assign mem[942 ] = 4'h0;
  assign mem[943 ] = 4'h4;
  assign mem[944 ] = 4'h0;
  assign mem[945 ] = 4'h1;
  assign mem[946 ] = 4'h0;
  assign mem[947 ] = 4'h2;
  assign mem[948 ] = 4'h0;
  assign mem[949 ] = 4'h1;
  assign mem[950 ] = 4'h0;
  assign mem[951 ] = 4'h3;
  assign mem[952 ] = 4'h0;
  assign mem[953 ] = 4'h1;
  assign mem[954 ] = 4'h0;
  assign mem[955 ] = 4'h2;
  assign mem[956 ] = 4'h0;
  assign mem[957 ] = 4'h1;
  assign mem[958 ] = 4'h0;
  assign mem[959 ] = 4'h6;
  assign mem[960 ] = 4'h0;
  assign mem[961 ] = 4'h1;
  assign mem[962 ] = 4'h0;
  assign mem[963 ] = 4'h2;
  assign mem[964 ] = 4'h0;
  assign mem[965 ] = 4'h1;
  assign mem[966 ] = 4'h0;
  assign mem[967 ] = 4'h3;
  assign mem[968 ] = 4'h0;
  assign mem[969 ] = 4'h1;
  assign mem[970 ] = 4'h0;
  assign mem[971 ] = 4'h2;
  assign mem[972 ] = 4'h0;
  assign mem[973 ] = 4'h1;
  assign mem[974 ] = 4'h0;
  assign mem[975 ] = 4'h4;
  assign mem[976 ] = 4'h0;
  assign mem[977 ] = 4'h1;
  assign mem[978 ] = 4'h0;
  assign mem[979 ] = 4'h2;
  assign mem[980 ] = 4'h0;
  assign mem[981 ] = 4'h1;
  assign mem[982 ] = 4'h0;
  assign mem[983 ] = 4'h3;
  assign mem[984 ] = 4'h0;
  assign mem[985 ] = 4'h1;
  assign mem[986 ] = 4'h0;
  assign mem[987 ] = 4'h2;
  assign mem[988 ] = 4'h0;
  assign mem[989 ] = 4'h1;
  assign mem[990 ] = 4'h0;
  assign mem[991 ] = 4'h5;
  assign mem[992 ] = 4'h0;
  assign mem[993 ] = 4'h1;
  assign mem[994 ] = 4'h0;
  assign mem[995 ] = 4'h2;
  assign mem[996 ] = 4'h0;
  assign mem[997 ] = 4'h1;
  assign mem[998 ] = 4'h0;
  assign mem[999 ] = 4'h3;
  assign mem[1000] = 4'h0;
  assign mem[1001] = 4'h1;
  assign mem[1002] = 4'h0;
  assign mem[1003] = 4'h2;
  assign mem[1004] = 4'h0;
  assign mem[1005] = 4'h1;
  assign mem[1006] = 4'h0;
  assign mem[1007] = 4'h4;
  assign mem[1008] = 4'h0;
  assign mem[1009] = 4'h1;
  assign mem[1010] = 4'h0;
  assign mem[1011] = 4'h2;
  assign mem[1012] = 4'h0;
  assign mem[1013] = 4'h1;
  assign mem[1014] = 4'h0;
  assign mem[1015] = 4'h3;
  assign mem[1016] = 4'h0;
  assign mem[1017] = 4'h1;
  assign mem[1018] = 4'h0;
  assign mem[1019] = 4'h2;
  assign mem[1020] = 4'h0;
  assign mem[1021] = 4'h1;
  assign mem[1022] = 4'h0;
  assign mem[1023] = 4'ha;
  assign mem[1024] = 4'h0;
  assign mem[1025] = 4'h1;
  assign mem[1026] = 4'h0;
  assign mem[1027] = 4'h2;
  assign mem[1028] = 4'h0;
  assign mem[1029] = 4'h1;
  assign mem[1030] = 4'h0;
  assign mem[1031] = 4'h3;
  assign mem[1032] = 4'h0;
  assign mem[1033] = 4'h1;
  assign mem[1034] = 4'h0;
  assign mem[1035] = 4'h2;
  assign mem[1036] = 4'h0;
  assign mem[1037] = 4'h1;
  assign mem[1038] = 4'h0;
  assign mem[1039] = 4'h4;
  assign mem[1040] = 4'h0;
  assign mem[1041] = 4'h1;
  assign mem[1042] = 4'h0;
  assign mem[1043] = 4'h2;
  assign mem[1044] = 4'h0;
  assign mem[1045] = 4'h1;
  assign mem[1046] = 4'h0;
  assign mem[1047] = 4'h3;
  assign mem[1048] = 4'h0;
  assign mem[1049] = 4'h1;
  assign mem[1050] = 4'h0;
  assign mem[1051] = 4'h2;
  assign mem[1052] = 4'h0;
  assign mem[1053] = 4'h1;
  assign mem[1054] = 4'h0;
  assign mem[1055] = 4'h5;
  assign mem[1056] = 4'h0;
  assign mem[1057] = 4'h1;
  assign mem[1058] = 4'h0;
  assign mem[1059] = 4'h2;
  assign mem[1060] = 4'h0;
  assign mem[1061] = 4'h1;
  assign mem[1062] = 4'h0;
  assign mem[1063] = 4'h3;
  assign mem[1064] = 4'h0;
  assign mem[1065] = 4'h1;
  assign mem[1066] = 4'h0;
  assign mem[1067] = 4'h2;
  assign mem[1068] = 4'h0;
  assign mem[1069] = 4'h1;
  assign mem[1070] = 4'h0;
  assign mem[1071] = 4'h4;
  assign mem[1072] = 4'h0;
  assign mem[1073] = 4'h1;
  assign mem[1074] = 4'h0;
  assign mem[1075] = 4'h2;
  assign mem[1076] = 4'h0;
  assign mem[1077] = 4'h1;
  assign mem[1078] = 4'h0;
  assign mem[1079] = 4'h3;
  assign mem[1080] = 4'h0;
  assign mem[1081] = 4'h1;
  assign mem[1082] = 4'h0;
  assign mem[1083] = 4'h2;
  assign mem[1084] = 4'h0;
  assign mem[1085] = 4'h1;
  assign mem[1086] = 4'h0;
  assign mem[1087] = 4'h6;
  assign mem[1088] = 4'h0;
  assign mem[1089] = 4'h1;
  assign mem[1090] = 4'h0;
  assign mem[1091] = 4'h2;
  assign mem[1092] = 4'h0;
  assign mem[1093] = 4'h1;
  assign mem[1094] = 4'h0;
  assign mem[1095] = 4'h3;
  assign mem[1096] = 4'h0;
  assign mem[1097] = 4'h1;
  assign mem[1098] = 4'h0;
  assign mem[1099] = 4'h2;
  assign mem[1100] = 4'h0;
  assign mem[1101] = 4'h1;
  assign mem[1102] = 4'h0;
  assign mem[1103] = 4'h4;
  assign mem[1104] = 4'h0;
  assign mem[1105] = 4'h1;
  assign mem[1106] = 4'h0;
  assign mem[1107] = 4'h2;
  assign mem[1108] = 4'h0;
  assign mem[1109] = 4'h1;
  assign mem[1110] = 4'h0;
  assign mem[1111] = 4'h3;
  assign mem[1112] = 4'h0;
  assign mem[1113] = 4'h1;
  assign mem[1114] = 4'h0;
  assign mem[1115] = 4'h2;
  assign mem[1116] = 4'h0;
  assign mem[1117] = 4'h1;
  assign mem[1118] = 4'h0;
  assign mem[1119] = 4'h5;
  assign mem[1120] = 4'h0;
  assign mem[1121] = 4'h1;
  assign mem[1122] = 4'h0;
  assign mem[1123] = 4'h2;
  assign mem[1124] = 4'h0;
  assign mem[1125] = 4'h1;
  assign mem[1126] = 4'h0;
  assign mem[1127] = 4'h3;
  assign mem[1128] = 4'h0;
  assign mem[1129] = 4'h1;
  assign mem[1130] = 4'h0;
  assign mem[1131] = 4'h2;
  assign mem[1132] = 4'h0;
  assign mem[1133] = 4'h1;
  assign mem[1134] = 4'h0;
  assign mem[1135] = 4'h4;
  assign mem[1136] = 4'h0;
  assign mem[1137] = 4'h1;
  assign mem[1138] = 4'h0;
  assign mem[1139] = 4'h2;
  assign mem[1140] = 4'h0;
  assign mem[1141] = 4'h1;
  assign mem[1142] = 4'h0;
  assign mem[1143] = 4'h3;
  assign mem[1144] = 4'h0;
  assign mem[1145] = 4'h1;
  assign mem[1146] = 4'h0;
  assign mem[1147] = 4'h2;
  assign mem[1148] = 4'h0;
  assign mem[1149] = 4'h1;
  assign mem[1150] = 4'h0;
  assign mem[1151] = 4'h7;
  assign mem[1152] = 4'h0;
  assign mem[1153] = 4'h1;
  assign mem[1154] = 4'h0;
  assign mem[1155] = 4'h2;
  assign mem[1156] = 4'h0;
  assign mem[1157] = 4'h1;
  assign mem[1158] = 4'h0;
  assign mem[1159] = 4'h3;
  assign mem[1160] = 4'h0;
  assign mem[1161] = 4'h1;
  assign mem[1162] = 4'h0;
  assign mem[1163] = 4'h2;
  assign mem[1164] = 4'h0;
  assign mem[1165] = 4'h1;
  assign mem[1166] = 4'h0;
  assign mem[1167] = 4'h4;
  assign mem[1168] = 4'h0;
  assign mem[1169] = 4'h1;
  assign mem[1170] = 4'h0;
  assign mem[1171] = 4'h2;
  assign mem[1172] = 4'h0;
  assign mem[1173] = 4'h1;
  assign mem[1174] = 4'h0;
  assign mem[1175] = 4'h3;
  assign mem[1176] = 4'h0;
  assign mem[1177] = 4'h1;
  assign mem[1178] = 4'h0;
  assign mem[1179] = 4'h2;
  assign mem[1180] = 4'h0;
  assign mem[1181] = 4'h1;
  assign mem[1182] = 4'h0;
  assign mem[1183] = 4'h5;
  assign mem[1184] = 4'h0;
  assign mem[1185] = 4'h1;
  assign mem[1186] = 4'h0;
  assign mem[1187] = 4'h2;
  assign mem[1188] = 4'h0;
  assign mem[1189] = 4'h1;
  assign mem[1190] = 4'h0;
  assign mem[1191] = 4'h3;
  assign mem[1192] = 4'h0;
  assign mem[1193] = 4'h1;
  assign mem[1194] = 4'h0;
  assign mem[1195] = 4'h2;
  assign mem[1196] = 4'h0;
  assign mem[1197] = 4'h1;
  assign mem[1198] = 4'h0;
  assign mem[1199] = 4'h4;
  assign mem[1200] = 4'h0;
  assign mem[1201] = 4'h1;
  assign mem[1202] = 4'h0;
  assign mem[1203] = 4'h2;
  assign mem[1204] = 4'h0;
  assign mem[1205] = 4'h1;
  assign mem[1206] = 4'h0;
  assign mem[1207] = 4'h3;
  assign mem[1208] = 4'h0;
  assign mem[1209] = 4'h1;
  assign mem[1210] = 4'h0;
  assign mem[1211] = 4'h2;
  assign mem[1212] = 4'h0;
  assign mem[1213] = 4'h1;
  assign mem[1214] = 4'h0;
  assign mem[1215] = 4'h6;
  assign mem[1216] = 4'h0;
  assign mem[1217] = 4'h1;
  assign mem[1218] = 4'h0;
  assign mem[1219] = 4'h2;
  assign mem[1220] = 4'h0;
  assign mem[1221] = 4'h1;
  assign mem[1222] = 4'h0;
  assign mem[1223] = 4'h3;
  assign mem[1224] = 4'h0;
  assign mem[1225] = 4'h1;
  assign mem[1226] = 4'h0;
  assign mem[1227] = 4'h2;
  assign mem[1228] = 4'h0;
  assign mem[1229] = 4'h1;
  assign mem[1230] = 4'h0;
  assign mem[1231] = 4'h4;
  assign mem[1232] = 4'h0;
  assign mem[1233] = 4'h1;
  assign mem[1234] = 4'h0;
  assign mem[1235] = 4'h2;
  assign mem[1236] = 4'h0;
  assign mem[1237] = 4'h1;
  assign mem[1238] = 4'h0;
  assign mem[1239] = 4'h3;
  assign mem[1240] = 4'h0;
  assign mem[1241] = 4'h1;
  assign mem[1242] = 4'h0;
  assign mem[1243] = 4'h2;
  assign mem[1244] = 4'h0;
  assign mem[1245] = 4'h1;
  assign mem[1246] = 4'h0;
  assign mem[1247] = 4'h5;
  assign mem[1248] = 4'h0;
  assign mem[1249] = 4'h1;
  assign mem[1250] = 4'h0;
  assign mem[1251] = 4'h2;
  assign mem[1252] = 4'h0;
  assign mem[1253] = 4'h1;
  assign mem[1254] = 4'h0;
  assign mem[1255] = 4'h3;
  assign mem[1256] = 4'h0;
  assign mem[1257] = 4'h1;
  assign mem[1258] = 4'h0;
  assign mem[1259] = 4'h2;
  assign mem[1260] = 4'h0;
  assign mem[1261] = 4'h1;
  assign mem[1262] = 4'h0;
  assign mem[1263] = 4'h4;
  assign mem[1264] = 4'h0;
  assign mem[1265] = 4'h1;
  assign mem[1266] = 4'h0;
  assign mem[1267] = 4'h2;
  assign mem[1268] = 4'h0;
  assign mem[1269] = 4'h1;
  assign mem[1270] = 4'h0;
  assign mem[1271] = 4'h3;
  assign mem[1272] = 4'h0;
  assign mem[1273] = 4'h1;
  assign mem[1274] = 4'h0;
  assign mem[1275] = 4'h2;
  assign mem[1276] = 4'h0;
  assign mem[1277] = 4'h1;
  assign mem[1278] = 4'h0;
  assign mem[1279] = 4'h8;
  assign mem[1280] = 4'h0;
  assign mem[1281] = 4'h1;
  assign mem[1282] = 4'h0;
  assign mem[1283] = 4'h2;
  assign mem[1284] = 4'h0;
  assign mem[1285] = 4'h1;
  assign mem[1286] = 4'h0;
  assign mem[1287] = 4'h3;
  assign mem[1288] = 4'h0;
  assign mem[1289] = 4'h1;
  assign mem[1290] = 4'h0;
  assign mem[1291] = 4'h2;
  assign mem[1292] = 4'h0;
  assign mem[1293] = 4'h1;
  assign mem[1294] = 4'h0;
  assign mem[1295] = 4'h4;
  assign mem[1296] = 4'h0;
  assign mem[1297] = 4'h1;
  assign mem[1298] = 4'h0;
  assign mem[1299] = 4'h2;
  assign mem[1300] = 4'h0;
  assign mem[1301] = 4'h1;
  assign mem[1302] = 4'h0;
  assign mem[1303] = 4'h3;
  assign mem[1304] = 4'h0;
  assign mem[1305] = 4'h1;
  assign mem[1306] = 4'h0;
  assign mem[1307] = 4'h2;
  assign mem[1308] = 4'h0;
  assign mem[1309] = 4'h1;
  assign mem[1310] = 4'h0;
  assign mem[1311] = 4'h5;
  assign mem[1312] = 4'h0;
  assign mem[1313] = 4'h1;
  assign mem[1314] = 4'h0;
  assign mem[1315] = 4'h2;
  assign mem[1316] = 4'h0;
  assign mem[1317] = 4'h1;
  assign mem[1318] = 4'h0;
  assign mem[1319] = 4'h3;
  assign mem[1320] = 4'h0;
  assign mem[1321] = 4'h1;
  assign mem[1322] = 4'h0;
  assign mem[1323] = 4'h2;
  assign mem[1324] = 4'h0;
  assign mem[1325] = 4'h1;
  assign mem[1326] = 4'h0;
  assign mem[1327] = 4'h4;
  assign mem[1328] = 4'h0;
  assign mem[1329] = 4'h1;
  assign mem[1330] = 4'h0;
  assign mem[1331] = 4'h2;
  assign mem[1332] = 4'h0;
  assign mem[1333] = 4'h1;
  assign mem[1334] = 4'h0;
  assign mem[1335] = 4'h3;
  assign mem[1336] = 4'h0;
  assign mem[1337] = 4'h1;
  assign mem[1338] = 4'h0;
  assign mem[1339] = 4'h2;
  assign mem[1340] = 4'h0;
  assign mem[1341] = 4'h1;
  assign mem[1342] = 4'h0;
  assign mem[1343] = 4'h6;
  assign mem[1344] = 4'h0;
  assign mem[1345] = 4'h1;
  assign mem[1346] = 4'h0;
  assign mem[1347] = 4'h2;
  assign mem[1348] = 4'h0;
  assign mem[1349] = 4'h1;
  assign mem[1350] = 4'h0;
  assign mem[1351] = 4'h3;
  assign mem[1352] = 4'h0;
  assign mem[1353] = 4'h1;
  assign mem[1354] = 4'h0;
  assign mem[1355] = 4'h2;
  assign mem[1356] = 4'h0;
  assign mem[1357] = 4'h1;
  assign mem[1358] = 4'h0;
  assign mem[1359] = 4'h4;
  assign mem[1360] = 4'h0;
  assign mem[1361] = 4'h1;
  assign mem[1362] = 4'h0;
  assign mem[1363] = 4'h2;
  assign mem[1364] = 4'h0;
  assign mem[1365] = 4'h1;
  assign mem[1366] = 4'h0;
  assign mem[1367] = 4'h3;
  assign mem[1368] = 4'h0;
  assign mem[1369] = 4'h1;
  assign mem[1370] = 4'h0;
  assign mem[1371] = 4'h2;
  assign mem[1372] = 4'h0;
  assign mem[1373] = 4'h1;
  assign mem[1374] = 4'h0;
  assign mem[1375] = 4'h5;
  assign mem[1376] = 4'h0;
  assign mem[1377] = 4'h1;
  assign mem[1378] = 4'h0;
  assign mem[1379] = 4'h2;
  assign mem[1380] = 4'h0;
  assign mem[1381] = 4'h1;
  assign mem[1382] = 4'h0;
  assign mem[1383] = 4'h3;
  assign mem[1384] = 4'h0;
  assign mem[1385] = 4'h1;
  assign mem[1386] = 4'h0;
  assign mem[1387] = 4'h2;
  assign mem[1388] = 4'h0;
  assign mem[1389] = 4'h1;
  assign mem[1390] = 4'h0;
  assign mem[1391] = 4'h4;
  assign mem[1392] = 4'h0;
  assign mem[1393] = 4'h1;
  assign mem[1394] = 4'h0;
  assign mem[1395] = 4'h2;
  assign mem[1396] = 4'h0;
  assign mem[1397] = 4'h1;
  assign mem[1398] = 4'h0;
  assign mem[1399] = 4'h3;
  assign mem[1400] = 4'h0;
  assign mem[1401] = 4'h1;
  assign mem[1402] = 4'h0;
  assign mem[1403] = 4'h2;
  assign mem[1404] = 4'h0;
  assign mem[1405] = 4'h1;
  assign mem[1406] = 4'h0;
  assign mem[1407] = 4'h7;
  assign mem[1408] = 4'h0;
  assign mem[1409] = 4'h1;
  assign mem[1410] = 4'h0;
  assign mem[1411] = 4'h2;
  assign mem[1412] = 4'h0;
  assign mem[1413] = 4'h1;
  assign mem[1414] = 4'h0;
  assign mem[1415] = 4'h3;
  assign mem[1416] = 4'h0;
  assign mem[1417] = 4'h1;
  assign mem[1418] = 4'h0;
  assign mem[1419] = 4'h2;
  assign mem[1420] = 4'h0;
  assign mem[1421] = 4'h1;
  assign mem[1422] = 4'h0;
  assign mem[1423] = 4'h4;
  assign mem[1424] = 4'h0;
  assign mem[1425] = 4'h1;
  assign mem[1426] = 4'h0;
  assign mem[1427] = 4'h2;
  assign mem[1428] = 4'h0;
  assign mem[1429] = 4'h1;
  assign mem[1430] = 4'h0;
  assign mem[1431] = 4'h3;
  assign mem[1432] = 4'h0;
  assign mem[1433] = 4'h1;
  assign mem[1434] = 4'h0;
  assign mem[1435] = 4'h2;
  assign mem[1436] = 4'h0;
  assign mem[1437] = 4'h1;
  assign mem[1438] = 4'h0;
  assign mem[1439] = 4'h5;
  assign mem[1440] = 4'h0;
  assign mem[1441] = 4'h1;
  assign mem[1442] = 4'h0;
  assign mem[1443] = 4'h2;
  assign mem[1444] = 4'h0;
  assign mem[1445] = 4'h1;
  assign mem[1446] = 4'h0;
  assign mem[1447] = 4'h3;
  assign mem[1448] = 4'h0;
  assign mem[1449] = 4'h1;
  assign mem[1450] = 4'h0;
  assign mem[1451] = 4'h2;
  assign mem[1452] = 4'h0;
  assign mem[1453] = 4'h1;
  assign mem[1454] = 4'h0;
  assign mem[1455] = 4'h4;
  assign mem[1456] = 4'h0;
  assign mem[1457] = 4'h1;
  assign mem[1458] = 4'h0;
  assign mem[1459] = 4'h2;
  assign mem[1460] = 4'h0;
  assign mem[1461] = 4'h1;
  assign mem[1462] = 4'h0;
  assign mem[1463] = 4'h3;
  assign mem[1464] = 4'h0;
  assign mem[1465] = 4'h1;
  assign mem[1466] = 4'h0;
  assign mem[1467] = 4'h2;
  assign mem[1468] = 4'h0;
  assign mem[1469] = 4'h1;
  assign mem[1470] = 4'h0;
  assign mem[1471] = 4'h6;
  assign mem[1472] = 4'h0;
  assign mem[1473] = 4'h1;
  assign mem[1474] = 4'h0;
  assign mem[1475] = 4'h2;
  assign mem[1476] = 4'h0;
  assign mem[1477] = 4'h1;
  assign mem[1478] = 4'h0;
  assign mem[1479] = 4'h3;
  assign mem[1480] = 4'h0;
  assign mem[1481] = 4'h1;
  assign mem[1482] = 4'h0;
  assign mem[1483] = 4'h2;
  assign mem[1484] = 4'h0;
  assign mem[1485] = 4'h1;
  assign mem[1486] = 4'h0;
  assign mem[1487] = 4'h4;
  assign mem[1488] = 4'h0;
  assign mem[1489] = 4'h1;
  assign mem[1490] = 4'h0;
  assign mem[1491] = 4'h2;
  assign mem[1492] = 4'h0;
  assign mem[1493] = 4'h1;
  assign mem[1494] = 4'h0;
  assign mem[1495] = 4'h3;
  assign mem[1496] = 4'h0;
  assign mem[1497] = 4'h1;
  assign mem[1498] = 4'h0;
  assign mem[1499] = 4'h2;
  assign mem[1500] = 4'h0;
  assign mem[1501] = 4'h1;
  assign mem[1502] = 4'h0;
  assign mem[1503] = 4'h5;
  assign mem[1504] = 4'h0;
  assign mem[1505] = 4'h1;
  assign mem[1506] = 4'h0;
  assign mem[1507] = 4'h2;
  assign mem[1508] = 4'h0;
  assign mem[1509] = 4'h1;
  assign mem[1510] = 4'h0;
  assign mem[1511] = 4'h3;
  assign mem[1512] = 4'h0;
  assign mem[1513] = 4'h1;
  assign mem[1514] = 4'h0;
  assign mem[1515] = 4'h2;
  assign mem[1516] = 4'h0;
  assign mem[1517] = 4'h1;
  assign mem[1518] = 4'h0;
  assign mem[1519] = 4'h4;
  assign mem[1520] = 4'h0;
  assign mem[1521] = 4'h1;
  assign mem[1522] = 4'h0;
  assign mem[1523] = 4'h2;
  assign mem[1524] = 4'h0;
  assign mem[1525] = 4'h1;
  assign mem[1526] = 4'h0;
  assign mem[1527] = 4'h3;
  assign mem[1528] = 4'h0;
  assign mem[1529] = 4'h1;
  assign mem[1530] = 4'h0;
  assign mem[1531] = 4'h2;
  assign mem[1532] = 4'h0;
  assign mem[1533] = 4'h1;
  assign mem[1534] = 4'h0;
  assign mem[1535] = 4'h9;
  assign mem[1536] = 4'h0;
  assign mem[1537] = 4'h1;
  assign mem[1538] = 4'h0;
  assign mem[1539] = 4'h2;
  assign mem[1540] = 4'h0;
  assign mem[1541] = 4'h1;
  assign mem[1542] = 4'h0;
  assign mem[1543] = 4'h3;
  assign mem[1544] = 4'h0;
  assign mem[1545] = 4'h1;
  assign mem[1546] = 4'h0;
  assign mem[1547] = 4'h2;
  assign mem[1548] = 4'h0;
  assign mem[1549] = 4'h1;
  assign mem[1550] = 4'h0;
  assign mem[1551] = 4'h4;
  assign mem[1552] = 4'h0;
  assign mem[1553] = 4'h1;
  assign mem[1554] = 4'h0;
  assign mem[1555] = 4'h2;
  assign mem[1556] = 4'h0;
  assign mem[1557] = 4'h1;
  assign mem[1558] = 4'h0;
  assign mem[1559] = 4'h3;
  assign mem[1560] = 4'h0;
  assign mem[1561] = 4'h1;
  assign mem[1562] = 4'h0;
  assign mem[1563] = 4'h2;
  assign mem[1564] = 4'h0;
  assign mem[1565] = 4'h1;
  assign mem[1566] = 4'h0;
  assign mem[1567] = 4'h5;
  assign mem[1568] = 4'h0;
  assign mem[1569] = 4'h1;
  assign mem[1570] = 4'h0;
  assign mem[1571] = 4'h2;
  assign mem[1572] = 4'h0;
  assign mem[1573] = 4'h1;
  assign mem[1574] = 4'h0;
  assign mem[1575] = 4'h3;
  assign mem[1576] = 4'h0;
  assign mem[1577] = 4'h1;
  assign mem[1578] = 4'h0;
  assign mem[1579] = 4'h2;
  assign mem[1580] = 4'h0;
  assign mem[1581] = 4'h1;
  assign mem[1582] = 4'h0;
  assign mem[1583] = 4'h4;
  assign mem[1584] = 4'h0;
  assign mem[1585] = 4'h1;
  assign mem[1586] = 4'h0;
  assign mem[1587] = 4'h2;
  assign mem[1588] = 4'h0;
  assign mem[1589] = 4'h1;
  assign mem[1590] = 4'h0;
  assign mem[1591] = 4'h3;
  assign mem[1592] = 4'h0;
  assign mem[1593] = 4'h1;
  assign mem[1594] = 4'h0;
  assign mem[1595] = 4'h2;
  assign mem[1596] = 4'h0;
  assign mem[1597] = 4'h1;
  assign mem[1598] = 4'h0;
  assign mem[1599] = 4'h6;
  assign mem[1600] = 4'h0;
  assign mem[1601] = 4'h1;
  assign mem[1602] = 4'h0;
  assign mem[1603] = 4'h2;
  assign mem[1604] = 4'h0;
  assign mem[1605] = 4'h1;
  assign mem[1606] = 4'h0;
  assign mem[1607] = 4'h3;
  assign mem[1608] = 4'h0;
  assign mem[1609] = 4'h1;
  assign mem[1610] = 4'h0;
  assign mem[1611] = 4'h2;
  assign mem[1612] = 4'h0;
  assign mem[1613] = 4'h1;
  assign mem[1614] = 4'h0;
  assign mem[1615] = 4'h4;
  assign mem[1616] = 4'h0;
  assign mem[1617] = 4'h1;
  assign mem[1618] = 4'h0;
  assign mem[1619] = 4'h2;
  assign mem[1620] = 4'h0;
  assign mem[1621] = 4'h1;
  assign mem[1622] = 4'h0;
  assign mem[1623] = 4'h3;
  assign mem[1624] = 4'h0;
  assign mem[1625] = 4'h1;
  assign mem[1626] = 4'h0;
  assign mem[1627] = 4'h2;
  assign mem[1628] = 4'h0;
  assign mem[1629] = 4'h1;
  assign mem[1630] = 4'h0;
  assign mem[1631] = 4'h5;
  assign mem[1632] = 4'h0;
  assign mem[1633] = 4'h1;
  assign mem[1634] = 4'h0;
  assign mem[1635] = 4'h2;
  assign mem[1636] = 4'h0;
  assign mem[1637] = 4'h1;
  assign mem[1638] = 4'h0;
  assign mem[1639] = 4'h3;
  assign mem[1640] = 4'h0;
  assign mem[1641] = 4'h1;
  assign mem[1642] = 4'h0;
  assign mem[1643] = 4'h2;
  assign mem[1644] = 4'h0;
  assign mem[1645] = 4'h1;
  assign mem[1646] = 4'h0;
  assign mem[1647] = 4'h4;
  assign mem[1648] = 4'h0;
  assign mem[1649] = 4'h1;
  assign mem[1650] = 4'h0;
  assign mem[1651] = 4'h2;
  assign mem[1652] = 4'h0;
  assign mem[1653] = 4'h1;
  assign mem[1654] = 4'h0;
  assign mem[1655] = 4'h3;
  assign mem[1656] = 4'h0;
  assign mem[1657] = 4'h1;
  assign mem[1658] = 4'h0;
  assign mem[1659] = 4'h2;
  assign mem[1660] = 4'h0;
  assign mem[1661] = 4'h1;
  assign mem[1662] = 4'h0;
  assign mem[1663] = 4'h7;
  assign mem[1664] = 4'h0;
  assign mem[1665] = 4'h1;
  assign mem[1666] = 4'h0;
  assign mem[1667] = 4'h2;
  assign mem[1668] = 4'h0;
  assign mem[1669] = 4'h1;
  assign mem[1670] = 4'h0;
  assign mem[1671] = 4'h3;
  assign mem[1672] = 4'h0;
  assign mem[1673] = 4'h1;
  assign mem[1674] = 4'h0;
  assign mem[1675] = 4'h2;
  assign mem[1676] = 4'h0;
  assign mem[1677] = 4'h1;
  assign mem[1678] = 4'h0;
  assign mem[1679] = 4'h4;
  assign mem[1680] = 4'h0;
  assign mem[1681] = 4'h1;
  assign mem[1682] = 4'h0;
  assign mem[1683] = 4'h2;
  assign mem[1684] = 4'h0;
  assign mem[1685] = 4'h1;
  assign mem[1686] = 4'h0;
  assign mem[1687] = 4'h3;
  assign mem[1688] = 4'h0;
  assign mem[1689] = 4'h1;
  assign mem[1690] = 4'h0;
  assign mem[1691] = 4'h2;
  assign mem[1692] = 4'h0;
  assign mem[1693] = 4'h1;
  assign mem[1694] = 4'h0;
  assign mem[1695] = 4'h5;
  assign mem[1696] = 4'h0;
  assign mem[1697] = 4'h1;
  assign mem[1698] = 4'h0;
  assign mem[1699] = 4'h2;
  assign mem[1700] = 4'h0;
  assign mem[1701] = 4'h1;
  assign mem[1702] = 4'h0;
  assign mem[1703] = 4'h3;
  assign mem[1704] = 4'h0;
  assign mem[1705] = 4'h1;
  assign mem[1706] = 4'h0;
  assign mem[1707] = 4'h2;
  assign mem[1708] = 4'h0;
  assign mem[1709] = 4'h1;
  assign mem[1710] = 4'h0;
  assign mem[1711] = 4'h4;
  assign mem[1712] = 4'h0;
  assign mem[1713] = 4'h1;
  assign mem[1714] = 4'h0;
  assign mem[1715] = 4'h2;
  assign mem[1716] = 4'h0;
  assign mem[1717] = 4'h1;
  assign mem[1718] = 4'h0;
  assign mem[1719] = 4'h3;
  assign mem[1720] = 4'h0;
  assign mem[1721] = 4'h1;
  assign mem[1722] = 4'h0;
  assign mem[1723] = 4'h2;
  assign mem[1724] = 4'h0;
  assign mem[1725] = 4'h1;
  assign mem[1726] = 4'h0;
  assign mem[1727] = 4'h6;
  assign mem[1728] = 4'h0;
  assign mem[1729] = 4'h1;
  assign mem[1730] = 4'h0;
  assign mem[1731] = 4'h2;
  assign mem[1732] = 4'h0;
  assign mem[1733] = 4'h1;
  assign mem[1734] = 4'h0;
  assign mem[1735] = 4'h3;
  assign mem[1736] = 4'h0;
  assign mem[1737] = 4'h1;
  assign mem[1738] = 4'h0;
  assign mem[1739] = 4'h2;
  assign mem[1740] = 4'h0;
  assign mem[1741] = 4'h1;
  assign mem[1742] = 4'h0;
  assign mem[1743] = 4'h4;
  assign mem[1744] = 4'h0;
  assign mem[1745] = 4'h1;
  assign mem[1746] = 4'h0;
  assign mem[1747] = 4'h2;
  assign mem[1748] = 4'h0;
  assign mem[1749] = 4'h1;
  assign mem[1750] = 4'h0;
  assign mem[1751] = 4'h3;
  assign mem[1752] = 4'h0;
  assign mem[1753] = 4'h1;
  assign mem[1754] = 4'h0;
  assign mem[1755] = 4'h2;
  assign mem[1756] = 4'h0;
  assign mem[1757] = 4'h1;
  assign mem[1758] = 4'h0;
  assign mem[1759] = 4'h5;
  assign mem[1760] = 4'h0;
  assign mem[1761] = 4'h1;
  assign mem[1762] = 4'h0;
  assign mem[1763] = 4'h2;
  assign mem[1764] = 4'h0;
  assign mem[1765] = 4'h1;
  assign mem[1766] = 4'h0;
  assign mem[1767] = 4'h3;
  assign mem[1768] = 4'h0;
  assign mem[1769] = 4'h1;
  assign mem[1770] = 4'h0;
  assign mem[1771] = 4'h2;
  assign mem[1772] = 4'h0;
  assign mem[1773] = 4'h1;
  assign mem[1774] = 4'h0;
  assign mem[1775] = 4'h4;
  assign mem[1776] = 4'h0;
  assign mem[1777] = 4'h1;
  assign mem[1778] = 4'h0;
  assign mem[1779] = 4'h2;
  assign mem[1780] = 4'h0;
  assign mem[1781] = 4'h1;
  assign mem[1782] = 4'h0;
  assign mem[1783] = 4'h3;
  assign mem[1784] = 4'h0;
  assign mem[1785] = 4'h1;
  assign mem[1786] = 4'h0;
  assign mem[1787] = 4'h2;
  assign mem[1788] = 4'h0;
  assign mem[1789] = 4'h1;
  assign mem[1790] = 4'h0;
  assign mem[1791] = 4'h8;
  assign mem[1792] = 4'h0;
  assign mem[1793] = 4'h1;
  assign mem[1794] = 4'h0;
  assign mem[1795] = 4'h2;
  assign mem[1796] = 4'h0;
  assign mem[1797] = 4'h1;
  assign mem[1798] = 4'h0;
  assign mem[1799] = 4'h3;
  assign mem[1800] = 4'h0;
  assign mem[1801] = 4'h1;
  assign mem[1802] = 4'h0;
  assign mem[1803] = 4'h2;
  assign mem[1804] = 4'h0;
  assign mem[1805] = 4'h1;
  assign mem[1806] = 4'h0;
  assign mem[1807] = 4'h4;
  assign mem[1808] = 4'h0;
  assign mem[1809] = 4'h1;
  assign mem[1810] = 4'h0;
  assign mem[1811] = 4'h2;
  assign mem[1812] = 4'h0;
  assign mem[1813] = 4'h1;
  assign mem[1814] = 4'h0;
  assign mem[1815] = 4'h3;
  assign mem[1816] = 4'h0;
  assign mem[1817] = 4'h1;
  assign mem[1818] = 4'h0;
  assign mem[1819] = 4'h2;
  assign mem[1820] = 4'h0;
  assign mem[1821] = 4'h1;
  assign mem[1822] = 4'h0;
  assign mem[1823] = 4'h5;
  assign mem[1824] = 4'h0;
  assign mem[1825] = 4'h1;
  assign mem[1826] = 4'h0;
  assign mem[1827] = 4'h2;
  assign mem[1828] = 4'h0;
  assign mem[1829] = 4'h1;
  assign mem[1830] = 4'h0;
  assign mem[1831] = 4'h3;
  assign mem[1832] = 4'h0;
  assign mem[1833] = 4'h1;
  assign mem[1834] = 4'h0;
  assign mem[1835] = 4'h2;
  assign mem[1836] = 4'h0;
  assign mem[1837] = 4'h1;
  assign mem[1838] = 4'h0;
  assign mem[1839] = 4'h4;
  assign mem[1840] = 4'h0;
  assign mem[1841] = 4'h1;
  assign mem[1842] = 4'h0;
  assign mem[1843] = 4'h2;
  assign mem[1844] = 4'h0;
  assign mem[1845] = 4'h1;
  assign mem[1846] = 4'h0;
  assign mem[1847] = 4'h3;
  assign mem[1848] = 4'h0;
  assign mem[1849] = 4'h1;
  assign mem[1850] = 4'h0;
  assign mem[1851] = 4'h2;
  assign mem[1852] = 4'h0;
  assign mem[1853] = 4'h1;
  assign mem[1854] = 4'h0;
  assign mem[1855] = 4'h6;
  assign mem[1856] = 4'h0;
  assign mem[1857] = 4'h1;
  assign mem[1858] = 4'h0;
  assign mem[1859] = 4'h2;
  assign mem[1860] = 4'h0;
  assign mem[1861] = 4'h1;
  assign mem[1862] = 4'h0;
  assign mem[1863] = 4'h3;
  assign mem[1864] = 4'h0;
  assign mem[1865] = 4'h1;
  assign mem[1866] = 4'h0;
  assign mem[1867] = 4'h2;
  assign mem[1868] = 4'h0;
  assign mem[1869] = 4'h1;
  assign mem[1870] = 4'h0;
  assign mem[1871] = 4'h4;
  assign mem[1872] = 4'h0;
  assign mem[1873] = 4'h1;
  assign mem[1874] = 4'h0;
  assign mem[1875] = 4'h2;
  assign mem[1876] = 4'h0;
  assign mem[1877] = 4'h1;
  assign mem[1878] = 4'h0;
  assign mem[1879] = 4'h3;
  assign mem[1880] = 4'h0;
  assign mem[1881] = 4'h1;
  assign mem[1882] = 4'h0;
  assign mem[1883] = 4'h2;
  assign mem[1884] = 4'h0;
  assign mem[1885] = 4'h1;
  assign mem[1886] = 4'h0;
  assign mem[1887] = 4'h5;
  assign mem[1888] = 4'h0;
  assign mem[1889] = 4'h1;
  assign mem[1890] = 4'h0;
  assign mem[1891] = 4'h2;
  assign mem[1892] = 4'h0;
  assign mem[1893] = 4'h1;
  assign mem[1894] = 4'h0;
  assign mem[1895] = 4'h3;
  assign mem[1896] = 4'h0;
  assign mem[1897] = 4'h1;
  assign mem[1898] = 4'h0;
  assign mem[1899] = 4'h2;
  assign mem[1900] = 4'h0;
  assign mem[1901] = 4'h1;
  assign mem[1902] = 4'h0;
  assign mem[1903] = 4'h4;
  assign mem[1904] = 4'h0;
  assign mem[1905] = 4'h1;
  assign mem[1906] = 4'h0;
  assign mem[1907] = 4'h2;
  assign mem[1908] = 4'h0;
  assign mem[1909] = 4'h1;
  assign mem[1910] = 4'h0;
  assign mem[1911] = 4'h3;
  assign mem[1912] = 4'h0;
  assign mem[1913] = 4'h1;
  assign mem[1914] = 4'h0;
  assign mem[1915] = 4'h2;
  assign mem[1916] = 4'h0;
  assign mem[1917] = 4'h1;
  assign mem[1918] = 4'h0;
  assign mem[1919] = 4'h7;
  assign mem[1920] = 4'h0;
  assign mem[1921] = 4'h1;
  assign mem[1922] = 4'h0;
  assign mem[1923] = 4'h2;
  assign mem[1924] = 4'h0;
  assign mem[1925] = 4'h1;
  assign mem[1926] = 4'h0;
  assign mem[1927] = 4'h3;
  assign mem[1928] = 4'h0;
  assign mem[1929] = 4'h1;
  assign mem[1930] = 4'h0;
  assign mem[1931] = 4'h2;
  assign mem[1932] = 4'h0;
  assign mem[1933] = 4'h1;
  assign mem[1934] = 4'h0;
  assign mem[1935] = 4'h4;
  assign mem[1936] = 4'h0;
  assign mem[1937] = 4'h1;
  assign mem[1938] = 4'h0;
  assign mem[1939] = 4'h2;
  assign mem[1940] = 4'h0;
  assign mem[1941] = 4'h1;
  assign mem[1942] = 4'h0;
  assign mem[1943] = 4'h3;
  assign mem[1944] = 4'h0;
  assign mem[1945] = 4'h1;
  assign mem[1946] = 4'h0;
  assign mem[1947] = 4'h2;
  assign mem[1948] = 4'h0;
  assign mem[1949] = 4'h1;
  assign mem[1950] = 4'h0;
  assign mem[1951] = 4'h5;
  assign mem[1952] = 4'h0;
  assign mem[1953] = 4'h1;
  assign mem[1954] = 4'h0;
  assign mem[1955] = 4'h2;
  assign mem[1956] = 4'h0;
  assign mem[1957] = 4'h1;
  assign mem[1958] = 4'h0;
  assign mem[1959] = 4'h3;
  assign mem[1960] = 4'h0;
  assign mem[1961] = 4'h1;
  assign mem[1962] = 4'h0;
  assign mem[1963] = 4'h2;
  assign mem[1964] = 4'h0;
  assign mem[1965] = 4'h1;
  assign mem[1966] = 4'h0;
  assign mem[1967] = 4'h4;
  assign mem[1968] = 4'h0;
  assign mem[1969] = 4'h1;
  assign mem[1970] = 4'h0;
  assign mem[1971] = 4'h2;
  assign mem[1972] = 4'h0;
  assign mem[1973] = 4'h1;
  assign mem[1974] = 4'h0;
  assign mem[1975] = 4'h3;
  assign mem[1976] = 4'h0;
  assign mem[1977] = 4'h1;
  assign mem[1978] = 4'h0;
  assign mem[1979] = 4'h2;
  assign mem[1980] = 4'h0;
  assign mem[1981] = 4'h1;
  assign mem[1982] = 4'h0;
  assign mem[1983] = 4'h6;
  assign mem[1984] = 4'h0;
  assign mem[1985] = 4'h1;
  assign mem[1986] = 4'h0;
  assign mem[1987] = 4'h2;
  assign mem[1988] = 4'h0;
  assign mem[1989] = 4'h1;
  assign mem[1990] = 4'h0;
  assign mem[1991] = 4'h3;
  assign mem[1992] = 4'h0;
  assign mem[1993] = 4'h1;
  assign mem[1994] = 4'h0;
  assign mem[1995] = 4'h2;
  assign mem[1996] = 4'h0;
  assign mem[1997] = 4'h1;
  assign mem[1998] = 4'h0;
  assign mem[1999] = 4'h4;
  assign mem[2000] = 4'h0;
  assign mem[2001] = 4'h1;
  assign mem[2002] = 4'h0;
  assign mem[2003] = 4'h2;
  assign mem[2004] = 4'h0;
  assign mem[2005] = 4'h1;
  assign mem[2006] = 4'h0;
  assign mem[2007] = 4'h3;
  assign mem[2008] = 4'h0;
  assign mem[2009] = 4'h1;
  assign mem[2010] = 4'h0;
  assign mem[2011] = 4'h2;
  assign mem[2012] = 4'h0;
  assign mem[2013] = 4'h1;
  assign mem[2014] = 4'h0;
  assign mem[2015] = 4'h5;
  assign mem[2016] = 4'h0;
  assign mem[2017] = 4'h1;
  assign mem[2018] = 4'h0;
  assign mem[2019] = 4'h2;
  assign mem[2020] = 4'h0;
  assign mem[2021] = 4'h1;
  assign mem[2022] = 4'h0;
  assign mem[2023] = 4'h3;
  assign mem[2024] = 4'h0;
  assign mem[2025] = 4'h1;
  assign mem[2026] = 4'h0;
  assign mem[2027] = 4'h2;
  assign mem[2028] = 4'h0;
  assign mem[2029] = 4'h1;
  assign mem[2030] = 4'h0;
  assign mem[2031] = 4'h4;
  assign mem[2032] = 4'h0;
  assign mem[2033] = 4'h1;
  assign mem[2034] = 4'h0;
  assign mem[2035] = 4'h2;
  assign mem[2036] = 4'h0;
  assign mem[2037] = 4'h1;
  assign mem[2038] = 4'h0;
  assign mem[2039] = 4'h3;
  assign mem[2040] = 4'h0;
  assign mem[2041] = 4'h1;
  assign mem[2042] = 4'h0;
  assign mem[2043] = 4'h2;
  assign mem[2044] = 4'h0;
  assign mem[2045] = 4'h1;
  assign mem[2046] = 4'h0;
  assign mem[2047] = 4'hb;
  assign mem[2048] = 4'h0;
  assign mem[2049] = 4'h1;
  assign mem[2050] = 4'h0;
  assign mem[2051] = 4'h2;
  assign mem[2052] = 4'h0;
  assign mem[2053] = 4'h1;
  assign mem[2054] = 4'h0;
  assign mem[2055] = 4'h3;
  assign mem[2056] = 4'h0;
  assign mem[2057] = 4'h1;
  assign mem[2058] = 4'h0;
  assign mem[2059] = 4'h2;
  assign mem[2060] = 4'h0;
  assign mem[2061] = 4'h1;
  assign mem[2062] = 4'h0;
  assign mem[2063] = 4'h4;
  assign mem[2064] = 4'h0;
  assign mem[2065] = 4'h1;
  assign mem[2066] = 4'h0;
  assign mem[2067] = 4'h2;
  assign mem[2068] = 4'h0;
  assign mem[2069] = 4'h1;
  assign mem[2070] = 4'h0;
  assign mem[2071] = 4'h3;
  assign mem[2072] = 4'h0;
  assign mem[2073] = 4'h1;
  assign mem[2074] = 4'h0;
  assign mem[2075] = 4'h2;
  assign mem[2076] = 4'h0;
  assign mem[2077] = 4'h1;
  assign mem[2078] = 4'h0;
  assign mem[2079] = 4'h5;
  assign mem[2080] = 4'h0;
  assign mem[2081] = 4'h1;
  assign mem[2082] = 4'h0;
  assign mem[2083] = 4'h2;
  assign mem[2084] = 4'h0;
  assign mem[2085] = 4'h1;
  assign mem[2086] = 4'h0;
  assign mem[2087] = 4'h3;
  assign mem[2088] = 4'h0;
  assign mem[2089] = 4'h1;
  assign mem[2090] = 4'h0;
  assign mem[2091] = 4'h2;
  assign mem[2092] = 4'h0;
  assign mem[2093] = 4'h1;
  assign mem[2094] = 4'h0;
  assign mem[2095] = 4'h4;
  assign mem[2096] = 4'h0;
  assign mem[2097] = 4'h1;
  assign mem[2098] = 4'h0;
  assign mem[2099] = 4'h2;
  assign mem[2100] = 4'h0;
  assign mem[2101] = 4'h1;
  assign mem[2102] = 4'h0;
  assign mem[2103] = 4'h3;
  assign mem[2104] = 4'h0;
  assign mem[2105] = 4'h1;
  assign mem[2106] = 4'h0;
  assign mem[2107] = 4'h2;
  assign mem[2108] = 4'h0;
  assign mem[2109] = 4'h1;
  assign mem[2110] = 4'h0;
  assign mem[2111] = 4'h6;
  assign mem[2112] = 4'h0;
  assign mem[2113] = 4'h1;
  assign mem[2114] = 4'h0;
  assign mem[2115] = 4'h2;
  assign mem[2116] = 4'h0;
  assign mem[2117] = 4'h1;
  assign mem[2118] = 4'h0;
  assign mem[2119] = 4'h3;
  assign mem[2120] = 4'h0;
  assign mem[2121] = 4'h1;
  assign mem[2122] = 4'h0;
  assign mem[2123] = 4'h2;
  assign mem[2124] = 4'h0;
  assign mem[2125] = 4'h1;
  assign mem[2126] = 4'h0;
  assign mem[2127] = 4'h4;
  assign mem[2128] = 4'h0;
  assign mem[2129] = 4'h1;
  assign mem[2130] = 4'h0;
  assign mem[2131] = 4'h2;
  assign mem[2132] = 4'h0;
  assign mem[2133] = 4'h1;
  assign mem[2134] = 4'h0;
  assign mem[2135] = 4'h3;
  assign mem[2136] = 4'h0;
  assign mem[2137] = 4'h1;
  assign mem[2138] = 4'h0;
  assign mem[2139] = 4'h2;
  assign mem[2140] = 4'h0;
  assign mem[2141] = 4'h1;
  assign mem[2142] = 4'h0;
  assign mem[2143] = 4'h5;
  assign mem[2144] = 4'h0;
  assign mem[2145] = 4'h1;
  assign mem[2146] = 4'h0;
  assign mem[2147] = 4'h2;
  assign mem[2148] = 4'h0;
  assign mem[2149] = 4'h1;
  assign mem[2150] = 4'h0;
  assign mem[2151] = 4'h3;
  assign mem[2152] = 4'h0;
  assign mem[2153] = 4'h1;
  assign mem[2154] = 4'h0;
  assign mem[2155] = 4'h2;
  assign mem[2156] = 4'h0;
  assign mem[2157] = 4'h1;
  assign mem[2158] = 4'h0;
  assign mem[2159] = 4'h4;
  assign mem[2160] = 4'h0;
  assign mem[2161] = 4'h1;
  assign mem[2162] = 4'h0;
  assign mem[2163] = 4'h2;
  assign mem[2164] = 4'h0;
  assign mem[2165] = 4'h1;
  assign mem[2166] = 4'h0;
  assign mem[2167] = 4'h3;
  assign mem[2168] = 4'h0;
  assign mem[2169] = 4'h1;
  assign mem[2170] = 4'h0;
  assign mem[2171] = 4'h2;
  assign mem[2172] = 4'h0;
  assign mem[2173] = 4'h1;
  assign mem[2174] = 4'h0;
  assign mem[2175] = 4'h7;
  assign mem[2176] = 4'h0;
  assign mem[2177] = 4'h1;
  assign mem[2178] = 4'h0;
  assign mem[2179] = 4'h2;
  assign mem[2180] = 4'h0;
  assign mem[2181] = 4'h1;
  assign mem[2182] = 4'h0;
  assign mem[2183] = 4'h3;
  assign mem[2184] = 4'h0;
  assign mem[2185] = 4'h1;
  assign mem[2186] = 4'h0;
  assign mem[2187] = 4'h2;
  assign mem[2188] = 4'h0;
  assign mem[2189] = 4'h1;
  assign mem[2190] = 4'h0;
  assign mem[2191] = 4'h4;
  assign mem[2192] = 4'h0;
  assign mem[2193] = 4'h1;
  assign mem[2194] = 4'h0;
  assign mem[2195] = 4'h2;
  assign mem[2196] = 4'h0;
  assign mem[2197] = 4'h1;
  assign mem[2198] = 4'h0;
  assign mem[2199] = 4'h3;
  assign mem[2200] = 4'h0;
  assign mem[2201] = 4'h1;
  assign mem[2202] = 4'h0;
  assign mem[2203] = 4'h2;
  assign mem[2204] = 4'h0;
  assign mem[2205] = 4'h1;
  assign mem[2206] = 4'h0;
  assign mem[2207] = 4'h5;
  assign mem[2208] = 4'h0;
  assign mem[2209] = 4'h1;
  assign mem[2210] = 4'h0;
  assign mem[2211] = 4'h2;
  assign mem[2212] = 4'h0;
  assign mem[2213] = 4'h1;
  assign mem[2214] = 4'h0;
  assign mem[2215] = 4'h3;
  assign mem[2216] = 4'h0;
  assign mem[2217] = 4'h1;
  assign mem[2218] = 4'h0;
  assign mem[2219] = 4'h2;
  assign mem[2220] = 4'h0;
  assign mem[2221] = 4'h1;
  assign mem[2222] = 4'h0;
  assign mem[2223] = 4'h4;
  assign mem[2224] = 4'h0;
  assign mem[2225] = 4'h1;
  assign mem[2226] = 4'h0;
  assign mem[2227] = 4'h2;
  assign mem[2228] = 4'h0;
  assign mem[2229] = 4'h1;
  assign mem[2230] = 4'h0;
  assign mem[2231] = 4'h3;
  assign mem[2232] = 4'h0;
  assign mem[2233] = 4'h1;
  assign mem[2234] = 4'h0;
  assign mem[2235] = 4'h2;
  assign mem[2236] = 4'h0;
  assign mem[2237] = 4'h1;
  assign mem[2238] = 4'h0;
  assign mem[2239] = 4'h6;
  assign mem[2240] = 4'h0;
  assign mem[2241] = 4'h1;
  assign mem[2242] = 4'h0;
  assign mem[2243] = 4'h2;
  assign mem[2244] = 4'h0;
  assign mem[2245] = 4'h1;
  assign mem[2246] = 4'h0;
  assign mem[2247] = 4'h3;
  assign mem[2248] = 4'h0;
  assign mem[2249] = 4'h1;
  assign mem[2250] = 4'h0;
  assign mem[2251] = 4'h2;
  assign mem[2252] = 4'h0;
  assign mem[2253] = 4'h1;
  assign mem[2254] = 4'h0;
  assign mem[2255] = 4'h4;
  assign mem[2256] = 4'h0;
  assign mem[2257] = 4'h1;
  assign mem[2258] = 4'h0;
  assign mem[2259] = 4'h2;
  assign mem[2260] = 4'h0;
  assign mem[2261] = 4'h1;
  assign mem[2262] = 4'h0;
  assign mem[2263] = 4'h3;
  assign mem[2264] = 4'h0;
  assign mem[2265] = 4'h1;
  assign mem[2266] = 4'h0;
  assign mem[2267] = 4'h2;
  assign mem[2268] = 4'h0;
  assign mem[2269] = 4'h1;
  assign mem[2270] = 4'h0;
  assign mem[2271] = 4'h5;
  assign mem[2272] = 4'h0;
  assign mem[2273] = 4'h1;
  assign mem[2274] = 4'h0;
  assign mem[2275] = 4'h2;
  assign mem[2276] = 4'h0;
  assign mem[2277] = 4'h1;
  assign mem[2278] = 4'h0;
  assign mem[2279] = 4'h3;
  assign mem[2280] = 4'h0;
  assign mem[2281] = 4'h1;
  assign mem[2282] = 4'h0;
  assign mem[2283] = 4'h2;
  assign mem[2284] = 4'h0;
  assign mem[2285] = 4'h1;
  assign mem[2286] = 4'h0;
  assign mem[2287] = 4'h4;
  assign mem[2288] = 4'h0;
  assign mem[2289] = 4'h1;
  assign mem[2290] = 4'h0;
  assign mem[2291] = 4'h2;
  assign mem[2292] = 4'h0;
  assign mem[2293] = 4'h1;
  assign mem[2294] = 4'h0;
  assign mem[2295] = 4'h3;
  assign mem[2296] = 4'h0;
  assign mem[2297] = 4'h1;
  assign mem[2298] = 4'h0;
  assign mem[2299] = 4'h2;
  assign mem[2300] = 4'h0;
  assign mem[2301] = 4'h1;
  assign mem[2302] = 4'h0;
  assign mem[2303] = 4'h8;
  assign mem[2304] = 4'h0;
  assign mem[2305] = 4'h1;
  assign mem[2306] = 4'h0;
  assign mem[2307] = 4'h2;
  assign mem[2308] = 4'h0;
  assign mem[2309] = 4'h1;
  assign mem[2310] = 4'h0;
  assign mem[2311] = 4'h3;
  assign mem[2312] = 4'h0;
  assign mem[2313] = 4'h1;
  assign mem[2314] = 4'h0;
  assign mem[2315] = 4'h2;
  assign mem[2316] = 4'h0;
  assign mem[2317] = 4'h1;
  assign mem[2318] = 4'h0;
  assign mem[2319] = 4'h4;
  assign mem[2320] = 4'h0;
  assign mem[2321] = 4'h1;
  assign mem[2322] = 4'h0;
  assign mem[2323] = 4'h2;
  assign mem[2324] = 4'h0;
  assign mem[2325] = 4'h1;
  assign mem[2326] = 4'h0;
  assign mem[2327] = 4'h3;
  assign mem[2328] = 4'h0;
  assign mem[2329] = 4'h1;
  assign mem[2330] = 4'h0;
  assign mem[2331] = 4'h2;
  assign mem[2332] = 4'h0;
  assign mem[2333] = 4'h1;
  assign mem[2334] = 4'h0;
  assign mem[2335] = 4'h5;
  assign mem[2336] = 4'h0;
  assign mem[2337] = 4'h1;
  assign mem[2338] = 4'h0;
  assign mem[2339] = 4'h2;
  assign mem[2340] = 4'h0;
  assign mem[2341] = 4'h1;
  assign mem[2342] = 4'h0;
  assign mem[2343] = 4'h3;
  assign mem[2344] = 4'h0;
  assign mem[2345] = 4'h1;
  assign mem[2346] = 4'h0;
  assign mem[2347] = 4'h2;
  assign mem[2348] = 4'h0;
  assign mem[2349] = 4'h1;
  assign mem[2350] = 4'h0;
  assign mem[2351] = 4'h4;
  assign mem[2352] = 4'h0;
  assign mem[2353] = 4'h1;
  assign mem[2354] = 4'h0;
  assign mem[2355] = 4'h2;
  assign mem[2356] = 4'h0;
  assign mem[2357] = 4'h1;
  assign mem[2358] = 4'h0;
  assign mem[2359] = 4'h3;
  assign mem[2360] = 4'h0;
  assign mem[2361] = 4'h1;
  assign mem[2362] = 4'h0;
  assign mem[2363] = 4'h2;
  assign mem[2364] = 4'h0;
  assign mem[2365] = 4'h1;
  assign mem[2366] = 4'h0;
  assign mem[2367] = 4'h6;
  assign mem[2368] = 4'h0;
  assign mem[2369] = 4'h1;
  assign mem[2370] = 4'h0;
  assign mem[2371] = 4'h2;
  assign mem[2372] = 4'h0;
  assign mem[2373] = 4'h1;
  assign mem[2374] = 4'h0;
  assign mem[2375] = 4'h3;
  assign mem[2376] = 4'h0;
  assign mem[2377] = 4'h1;
  assign mem[2378] = 4'h0;
  assign mem[2379] = 4'h2;
  assign mem[2380] = 4'h0;
  assign mem[2381] = 4'h1;
  assign mem[2382] = 4'h0;
  assign mem[2383] = 4'h4;
  assign mem[2384] = 4'h0;
  assign mem[2385] = 4'h1;
  assign mem[2386] = 4'h0;
  assign mem[2387] = 4'h2;
  assign mem[2388] = 4'h0;
  assign mem[2389] = 4'h1;
  assign mem[2390] = 4'h0;
  assign mem[2391] = 4'h3;
  assign mem[2392] = 4'h0;
  assign mem[2393] = 4'h1;
  assign mem[2394] = 4'h0;
  assign mem[2395] = 4'h2;
  assign mem[2396] = 4'h0;
  assign mem[2397] = 4'h1;
  assign mem[2398] = 4'h0;
  assign mem[2399] = 4'h5;
  assign mem[2400] = 4'h0;
  assign mem[2401] = 4'h1;
  assign mem[2402] = 4'h0;
  assign mem[2403] = 4'h2;
  assign mem[2404] = 4'h0;
  assign mem[2405] = 4'h1;
  assign mem[2406] = 4'h0;
  assign mem[2407] = 4'h3;
  assign mem[2408] = 4'h0;
  assign mem[2409] = 4'h1;
  assign mem[2410] = 4'h0;
  assign mem[2411] = 4'h2;
  assign mem[2412] = 4'h0;
  assign mem[2413] = 4'h1;
  assign mem[2414] = 4'h0;
  assign mem[2415] = 4'h4;
  assign mem[2416] = 4'h0;
  assign mem[2417] = 4'h1;
  assign mem[2418] = 4'h0;
  assign mem[2419] = 4'h2;
  assign mem[2420] = 4'h0;
  assign mem[2421] = 4'h1;
  assign mem[2422] = 4'h0;
  assign mem[2423] = 4'h3;
  assign mem[2424] = 4'h0;
  assign mem[2425] = 4'h1;
  assign mem[2426] = 4'h0;
  assign mem[2427] = 4'h2;
  assign mem[2428] = 4'h0;
  assign mem[2429] = 4'h1;
  assign mem[2430] = 4'h0;
  assign mem[2431] = 4'h7;
  assign mem[2432] = 4'h0;
  assign mem[2433] = 4'h1;
  assign mem[2434] = 4'h0;
  assign mem[2435] = 4'h2;
  assign mem[2436] = 4'h0;
  assign mem[2437] = 4'h1;
  assign mem[2438] = 4'h0;
  assign mem[2439] = 4'h3;
  assign mem[2440] = 4'h0;
  assign mem[2441] = 4'h1;
  assign mem[2442] = 4'h0;
  assign mem[2443] = 4'h2;
  assign mem[2444] = 4'h0;
  assign mem[2445] = 4'h1;
  assign mem[2446] = 4'h0;
  assign mem[2447] = 4'h4;
  assign mem[2448] = 4'h0;
  assign mem[2449] = 4'h1;
  assign mem[2450] = 4'h0;
  assign mem[2451] = 4'h2;
  assign mem[2452] = 4'h0;
  assign mem[2453] = 4'h1;
  assign mem[2454] = 4'h0;
  assign mem[2455] = 4'h3;
  assign mem[2456] = 4'h0;
  assign mem[2457] = 4'h1;
  assign mem[2458] = 4'h0;
  assign mem[2459] = 4'h2;
  assign mem[2460] = 4'h0;
  assign mem[2461] = 4'h1;
  assign mem[2462] = 4'h0;
  assign mem[2463] = 4'h5;
  assign mem[2464] = 4'h0;
  assign mem[2465] = 4'h1;
  assign mem[2466] = 4'h0;
  assign mem[2467] = 4'h2;
  assign mem[2468] = 4'h0;
  assign mem[2469] = 4'h1;
  assign mem[2470] = 4'h0;
  assign mem[2471] = 4'h3;
  assign mem[2472] = 4'h0;
  assign mem[2473] = 4'h1;
  assign mem[2474] = 4'h0;
  assign mem[2475] = 4'h2;
  assign mem[2476] = 4'h0;
  assign mem[2477] = 4'h1;
  assign mem[2478] = 4'h0;
  assign mem[2479] = 4'h4;
  assign mem[2480] = 4'h0;
  assign mem[2481] = 4'h1;
  assign mem[2482] = 4'h0;
  assign mem[2483] = 4'h2;
  assign mem[2484] = 4'h0;
  assign mem[2485] = 4'h1;
  assign mem[2486] = 4'h0;
  assign mem[2487] = 4'h3;
  assign mem[2488] = 4'h0;
  assign mem[2489] = 4'h1;
  assign mem[2490] = 4'h0;
  assign mem[2491] = 4'h2;
  assign mem[2492] = 4'h0;
  assign mem[2493] = 4'h1;
  assign mem[2494] = 4'h0;
  assign mem[2495] = 4'h6;
  assign mem[2496] = 4'h0;
  assign mem[2497] = 4'h1;
  assign mem[2498] = 4'h0;
  assign mem[2499] = 4'h2;
  assign mem[2500] = 4'h0;
  assign mem[2501] = 4'h1;
  assign mem[2502] = 4'h0;
  assign mem[2503] = 4'h3;
  assign mem[2504] = 4'h0;
  assign mem[2505] = 4'h1;
  assign mem[2506] = 4'h0;
  assign mem[2507] = 4'h2;
  assign mem[2508] = 4'h0;
  assign mem[2509] = 4'h1;
  assign mem[2510] = 4'h0;
  assign mem[2511] = 4'h4;
  assign mem[2512] = 4'h0;
  assign mem[2513] = 4'h1;
  assign mem[2514] = 4'h0;
  assign mem[2515] = 4'h2;
  assign mem[2516] = 4'h0;
  assign mem[2517] = 4'h1;
  assign mem[2518] = 4'h0;
  assign mem[2519] = 4'h3;
  assign mem[2520] = 4'h0;
  assign mem[2521] = 4'h1;
  assign mem[2522] = 4'h0;
  assign mem[2523] = 4'h2;
  assign mem[2524] = 4'h0;
  assign mem[2525] = 4'h1;
  assign mem[2526] = 4'h0;
  assign mem[2527] = 4'h5;
  assign mem[2528] = 4'h0;
  assign mem[2529] = 4'h1;
  assign mem[2530] = 4'h0;
  assign mem[2531] = 4'h2;
  assign mem[2532] = 4'h0;
  assign mem[2533] = 4'h1;
  assign mem[2534] = 4'h0;
  assign mem[2535] = 4'h3;
  assign mem[2536] = 4'h0;
  assign mem[2537] = 4'h1;
  assign mem[2538] = 4'h0;
  assign mem[2539] = 4'h2;
  assign mem[2540] = 4'h0;
  assign mem[2541] = 4'h1;
  assign mem[2542] = 4'h0;
  assign mem[2543] = 4'h4;
  assign mem[2544] = 4'h0;
  assign mem[2545] = 4'h1;
  assign mem[2546] = 4'h0;
  assign mem[2547] = 4'h2;
  assign mem[2548] = 4'h0;
  assign mem[2549] = 4'h1;
  assign mem[2550] = 4'h0;
  assign mem[2551] = 4'h3;
  assign mem[2552] = 4'h0;
  assign mem[2553] = 4'h1;
  assign mem[2554] = 4'h0;
  assign mem[2555] = 4'h2;
  assign mem[2556] = 4'h0;
  assign mem[2557] = 4'h1;
  assign mem[2558] = 4'h0;
  assign mem[2559] = 4'h9;
  assign mem[2560] = 4'h0;
  assign mem[2561] = 4'h1;
  assign mem[2562] = 4'h0;
  assign mem[2563] = 4'h2;
  assign mem[2564] = 4'h0;
  assign mem[2565] = 4'h1;
  assign mem[2566] = 4'h0;
  assign mem[2567] = 4'h3;
  assign mem[2568] = 4'h0;
  assign mem[2569] = 4'h1;
  assign mem[2570] = 4'h0;
  assign mem[2571] = 4'h2;
  assign mem[2572] = 4'h0;
  assign mem[2573] = 4'h1;
  assign mem[2574] = 4'h0;
  assign mem[2575] = 4'h4;
  assign mem[2576] = 4'h0;
  assign mem[2577] = 4'h1;
  assign mem[2578] = 4'h0;
  assign mem[2579] = 4'h2;
  assign mem[2580] = 4'h0;
  assign mem[2581] = 4'h1;
  assign mem[2582] = 4'h0;
  assign mem[2583] = 4'h3;
  assign mem[2584] = 4'h0;
  assign mem[2585] = 4'h1;
  assign mem[2586] = 4'h0;
  assign mem[2587] = 4'h2;
  assign mem[2588] = 4'h0;
  assign mem[2589] = 4'h1;
  assign mem[2590] = 4'h0;
  assign mem[2591] = 4'h5;
  assign mem[2592] = 4'h0;
  assign mem[2593] = 4'h1;
  assign mem[2594] = 4'h0;
  assign mem[2595] = 4'h2;
  assign mem[2596] = 4'h0;
  assign mem[2597] = 4'h1;
  assign mem[2598] = 4'h0;
  assign mem[2599] = 4'h3;
  assign mem[2600] = 4'h0;
  assign mem[2601] = 4'h1;
  assign mem[2602] = 4'h0;
  assign mem[2603] = 4'h2;
  assign mem[2604] = 4'h0;
  assign mem[2605] = 4'h1;
  assign mem[2606] = 4'h0;
  assign mem[2607] = 4'h4;
  assign mem[2608] = 4'h0;
  assign mem[2609] = 4'h1;
  assign mem[2610] = 4'h0;
  assign mem[2611] = 4'h2;
  assign mem[2612] = 4'h0;
  assign mem[2613] = 4'h1;
  assign mem[2614] = 4'h0;
  assign mem[2615] = 4'h3;
  assign mem[2616] = 4'h0;
  assign mem[2617] = 4'h1;
  assign mem[2618] = 4'h0;
  assign mem[2619] = 4'h2;
  assign mem[2620] = 4'h0;
  assign mem[2621] = 4'h1;
  assign mem[2622] = 4'h0;
  assign mem[2623] = 4'h6;
  assign mem[2624] = 4'h0;
  assign mem[2625] = 4'h1;
  assign mem[2626] = 4'h0;
  assign mem[2627] = 4'h2;
  assign mem[2628] = 4'h0;
  assign mem[2629] = 4'h1;
  assign mem[2630] = 4'h0;
  assign mem[2631] = 4'h3;
  assign mem[2632] = 4'h0;
  assign mem[2633] = 4'h1;
  assign mem[2634] = 4'h0;
  assign mem[2635] = 4'h2;
  assign mem[2636] = 4'h0;
  assign mem[2637] = 4'h1;
  assign mem[2638] = 4'h0;
  assign mem[2639] = 4'h4;
  assign mem[2640] = 4'h0;
  assign mem[2641] = 4'h1;
  assign mem[2642] = 4'h0;
  assign mem[2643] = 4'h2;
  assign mem[2644] = 4'h0;
  assign mem[2645] = 4'h1;
  assign mem[2646] = 4'h0;
  assign mem[2647] = 4'h3;
  assign mem[2648] = 4'h0;
  assign mem[2649] = 4'h1;
  assign mem[2650] = 4'h0;
  assign mem[2651] = 4'h2;
  assign mem[2652] = 4'h0;
  assign mem[2653] = 4'h1;
  assign mem[2654] = 4'h0;
  assign mem[2655] = 4'h5;
  assign mem[2656] = 4'h0;
  assign mem[2657] = 4'h1;
  assign mem[2658] = 4'h0;
  assign mem[2659] = 4'h2;
  assign mem[2660] = 4'h0;
  assign mem[2661] = 4'h1;
  assign mem[2662] = 4'h0;
  assign mem[2663] = 4'h3;
  assign mem[2664] = 4'h0;
  assign mem[2665] = 4'h1;
  assign mem[2666] = 4'h0;
  assign mem[2667] = 4'h2;
  assign mem[2668] = 4'h0;
  assign mem[2669] = 4'h1;
  assign mem[2670] = 4'h0;
  assign mem[2671] = 4'h4;
  assign mem[2672] = 4'h0;
  assign mem[2673] = 4'h1;
  assign mem[2674] = 4'h0;
  assign mem[2675] = 4'h2;
  assign mem[2676] = 4'h0;
  assign mem[2677] = 4'h1;
  assign mem[2678] = 4'h0;
  assign mem[2679] = 4'h3;
  assign mem[2680] = 4'h0;
  assign mem[2681] = 4'h1;
  assign mem[2682] = 4'h0;
  assign mem[2683] = 4'h2;
  assign mem[2684] = 4'h0;
  assign mem[2685] = 4'h1;
  assign mem[2686] = 4'h0;
  assign mem[2687] = 4'h7;
  assign mem[2688] = 4'h0;
  assign mem[2689] = 4'h1;
  assign mem[2690] = 4'h0;
  assign mem[2691] = 4'h2;
  assign mem[2692] = 4'h0;
  assign mem[2693] = 4'h1;
  assign mem[2694] = 4'h0;
  assign mem[2695] = 4'h3;
  assign mem[2696] = 4'h0;
  assign mem[2697] = 4'h1;
  assign mem[2698] = 4'h0;
  assign mem[2699] = 4'h2;
  assign mem[2700] = 4'h0;
  assign mem[2701] = 4'h1;
  assign mem[2702] = 4'h0;
  assign mem[2703] = 4'h4;
  assign mem[2704] = 4'h0;
  assign mem[2705] = 4'h1;
  assign mem[2706] = 4'h0;
  assign mem[2707] = 4'h2;
  assign mem[2708] = 4'h0;
  assign mem[2709] = 4'h1;
  assign mem[2710] = 4'h0;
  assign mem[2711] = 4'h3;
  assign mem[2712] = 4'h0;
  assign mem[2713] = 4'h1;
  assign mem[2714] = 4'h0;
  assign mem[2715] = 4'h2;
  assign mem[2716] = 4'h0;
  assign mem[2717] = 4'h1;
  assign mem[2718] = 4'h0;
  assign mem[2719] = 4'h5;
  assign mem[2720] = 4'h0;
  assign mem[2721] = 4'h1;
  assign mem[2722] = 4'h0;
  assign mem[2723] = 4'h2;
  assign mem[2724] = 4'h0;
  assign mem[2725] = 4'h1;
  assign mem[2726] = 4'h0;
  assign mem[2727] = 4'h3;
  assign mem[2728] = 4'h0;
  assign mem[2729] = 4'h1;
  assign mem[2730] = 4'h0;
  assign mem[2731] = 4'h2;
  assign mem[2732] = 4'h0;
  assign mem[2733] = 4'h1;
  assign mem[2734] = 4'h0;
  assign mem[2735] = 4'h4;
  assign mem[2736] = 4'h0;
  assign mem[2737] = 4'h1;
  assign mem[2738] = 4'h0;
  assign mem[2739] = 4'h2;
  assign mem[2740] = 4'h0;
  assign mem[2741] = 4'h1;
  assign mem[2742] = 4'h0;
  assign mem[2743] = 4'h3;
  assign mem[2744] = 4'h0;
  assign mem[2745] = 4'h1;
  assign mem[2746] = 4'h0;
  assign mem[2747] = 4'h2;
  assign mem[2748] = 4'h0;
  assign mem[2749] = 4'h1;
  assign mem[2750] = 4'h0;
  assign mem[2751] = 4'h6;
  assign mem[2752] = 4'h0;
  assign mem[2753] = 4'h1;
  assign mem[2754] = 4'h0;
  assign mem[2755] = 4'h2;
  assign mem[2756] = 4'h0;
  assign mem[2757] = 4'h1;
  assign mem[2758] = 4'h0;
  assign mem[2759] = 4'h3;
  assign mem[2760] = 4'h0;
  assign mem[2761] = 4'h1;
  assign mem[2762] = 4'h0;
  assign mem[2763] = 4'h2;
  assign mem[2764] = 4'h0;
  assign mem[2765] = 4'h1;
  assign mem[2766] = 4'h0;
  assign mem[2767] = 4'h4;
  assign mem[2768] = 4'h0;
  assign mem[2769] = 4'h1;
  assign mem[2770] = 4'h0;
  assign mem[2771] = 4'h2;
  assign mem[2772] = 4'h0;
  assign mem[2773] = 4'h1;
  assign mem[2774] = 4'h0;
  assign mem[2775] = 4'h3;
  assign mem[2776] = 4'h0;
  assign mem[2777] = 4'h1;
  assign mem[2778] = 4'h0;
  assign mem[2779] = 4'h2;
  assign mem[2780] = 4'h0;
  assign mem[2781] = 4'h1;
  assign mem[2782] = 4'h0;
  assign mem[2783] = 4'h5;
  assign mem[2784] = 4'h0;
  assign mem[2785] = 4'h1;
  assign mem[2786] = 4'h0;
  assign mem[2787] = 4'h2;
  assign mem[2788] = 4'h0;
  assign mem[2789] = 4'h1;
  assign mem[2790] = 4'h0;
  assign mem[2791] = 4'h3;
  assign mem[2792] = 4'h0;
  assign mem[2793] = 4'h1;
  assign mem[2794] = 4'h0;
  assign mem[2795] = 4'h2;
  assign mem[2796] = 4'h0;
  assign mem[2797] = 4'h1;
  assign mem[2798] = 4'h0;
  assign mem[2799] = 4'h4;
  assign mem[2800] = 4'h0;
  assign mem[2801] = 4'h1;
  assign mem[2802] = 4'h0;
  assign mem[2803] = 4'h2;
  assign mem[2804] = 4'h0;
  assign mem[2805] = 4'h1;
  assign mem[2806] = 4'h0;
  assign mem[2807] = 4'h3;
  assign mem[2808] = 4'h0;
  assign mem[2809] = 4'h1;
  assign mem[2810] = 4'h0;
  assign mem[2811] = 4'h2;
  assign mem[2812] = 4'h0;
  assign mem[2813] = 4'h1;
  assign mem[2814] = 4'h0;
  assign mem[2815] = 4'h8;
  assign mem[2816] = 4'h0;
  assign mem[2817] = 4'h1;
  assign mem[2818] = 4'h0;
  assign mem[2819] = 4'h2;
  assign mem[2820] = 4'h0;
  assign mem[2821] = 4'h1;
  assign mem[2822] = 4'h0;
  assign mem[2823] = 4'h3;
  assign mem[2824] = 4'h0;
  assign mem[2825] = 4'h1;
  assign mem[2826] = 4'h0;
  assign mem[2827] = 4'h2;
  assign mem[2828] = 4'h0;
  assign mem[2829] = 4'h1;
  assign mem[2830] = 4'h0;
  assign mem[2831] = 4'h4;
  assign mem[2832] = 4'h0;
  assign mem[2833] = 4'h1;
  assign mem[2834] = 4'h0;
  assign mem[2835] = 4'h2;
  assign mem[2836] = 4'h0;
  assign mem[2837] = 4'h1;
  assign mem[2838] = 4'h0;
  assign mem[2839] = 4'h3;
  assign mem[2840] = 4'h0;
  assign mem[2841] = 4'h1;
  assign mem[2842] = 4'h0;
  assign mem[2843] = 4'h2;
  assign mem[2844] = 4'h0;
  assign mem[2845] = 4'h1;
  assign mem[2846] = 4'h0;
  assign mem[2847] = 4'h5;
  assign mem[2848] = 4'h0;
  assign mem[2849] = 4'h1;
  assign mem[2850] = 4'h0;
  assign mem[2851] = 4'h2;
  assign mem[2852] = 4'h0;
  assign mem[2853] = 4'h1;
  assign mem[2854] = 4'h0;
  assign mem[2855] = 4'h3;
  assign mem[2856] = 4'h0;
  assign mem[2857] = 4'h1;
  assign mem[2858] = 4'h0;
  assign mem[2859] = 4'h2;
  assign mem[2860] = 4'h0;
  assign mem[2861] = 4'h1;
  assign mem[2862] = 4'h0;
  assign mem[2863] = 4'h4;
  assign mem[2864] = 4'h0;
  assign mem[2865] = 4'h1;
  assign mem[2866] = 4'h0;
  assign mem[2867] = 4'h2;
  assign mem[2868] = 4'h0;
  assign mem[2869] = 4'h1;
  assign mem[2870] = 4'h0;
  assign mem[2871] = 4'h3;
  assign mem[2872] = 4'h0;
  assign mem[2873] = 4'h1;
  assign mem[2874] = 4'h0;
  assign mem[2875] = 4'h2;
  assign mem[2876] = 4'h0;
  assign mem[2877] = 4'h1;
  assign mem[2878] = 4'h0;
  assign mem[2879] = 4'h6;
  assign mem[2880] = 4'h0;
  assign mem[2881] = 4'h1;
  assign mem[2882] = 4'h0;
  assign mem[2883] = 4'h2;
  assign mem[2884] = 4'h0;
  assign mem[2885] = 4'h1;
  assign mem[2886] = 4'h0;
  assign mem[2887] = 4'h3;
  assign mem[2888] = 4'h0;
  assign mem[2889] = 4'h1;
  assign mem[2890] = 4'h0;
  assign mem[2891] = 4'h2;
  assign mem[2892] = 4'h0;
  assign mem[2893] = 4'h1;
  assign mem[2894] = 4'h0;
  assign mem[2895] = 4'h4;
  assign mem[2896] = 4'h0;
  assign mem[2897] = 4'h1;
  assign mem[2898] = 4'h0;
  assign mem[2899] = 4'h2;
  assign mem[2900] = 4'h0;
  assign mem[2901] = 4'h1;
  assign mem[2902] = 4'h0;
  assign mem[2903] = 4'h3;
  assign mem[2904] = 4'h0;
  assign mem[2905] = 4'h1;
  assign mem[2906] = 4'h0;
  assign mem[2907] = 4'h2;
  assign mem[2908] = 4'h0;
  assign mem[2909] = 4'h1;
  assign mem[2910] = 4'h0;
  assign mem[2911] = 4'h5;
  assign mem[2912] = 4'h0;
  assign mem[2913] = 4'h1;
  assign mem[2914] = 4'h0;
  assign mem[2915] = 4'h2;
  assign mem[2916] = 4'h0;
  assign mem[2917] = 4'h1;
  assign mem[2918] = 4'h0;
  assign mem[2919] = 4'h3;
  assign mem[2920] = 4'h0;
  assign mem[2921] = 4'h1;
  assign mem[2922] = 4'h0;
  assign mem[2923] = 4'h2;
  assign mem[2924] = 4'h0;
  assign mem[2925] = 4'h1;
  assign mem[2926] = 4'h0;
  assign mem[2927] = 4'h4;
  assign mem[2928] = 4'h0;
  assign mem[2929] = 4'h1;
  assign mem[2930] = 4'h0;
  assign mem[2931] = 4'h2;
  assign mem[2932] = 4'h0;
  assign mem[2933] = 4'h1;
  assign mem[2934] = 4'h0;
  assign mem[2935] = 4'h3;
  assign mem[2936] = 4'h0;
  assign mem[2937] = 4'h1;
  assign mem[2938] = 4'h0;
  assign mem[2939] = 4'h2;
  assign mem[2940] = 4'h0;
  assign mem[2941] = 4'h1;
  assign mem[2942] = 4'h0;
  assign mem[2943] = 4'h7;
  assign mem[2944] = 4'h0;
  assign mem[2945] = 4'h1;
  assign mem[2946] = 4'h0;
  assign mem[2947] = 4'h2;
  assign mem[2948] = 4'h0;
  assign mem[2949] = 4'h1;
  assign mem[2950] = 4'h0;
  assign mem[2951] = 4'h3;
  assign mem[2952] = 4'h0;
  assign mem[2953] = 4'h1;
  assign mem[2954] = 4'h0;
  assign mem[2955] = 4'h2;
  assign mem[2956] = 4'h0;
  assign mem[2957] = 4'h1;
  assign mem[2958] = 4'h0;
  assign mem[2959] = 4'h4;
  assign mem[2960] = 4'h0;
  assign mem[2961] = 4'h1;
  assign mem[2962] = 4'h0;
  assign mem[2963] = 4'h2;
  assign mem[2964] = 4'h0;
  assign mem[2965] = 4'h1;
  assign mem[2966] = 4'h0;
  assign mem[2967] = 4'h3;
  assign mem[2968] = 4'h0;
  assign mem[2969] = 4'h1;
  assign mem[2970] = 4'h0;
  assign mem[2971] = 4'h2;
  assign mem[2972] = 4'h0;
  assign mem[2973] = 4'h1;
  assign mem[2974] = 4'h0;
  assign mem[2975] = 4'h5;
  assign mem[2976] = 4'h0;
  assign mem[2977] = 4'h1;
  assign mem[2978] = 4'h0;
  assign mem[2979] = 4'h2;
  assign mem[2980] = 4'h0;
  assign mem[2981] = 4'h1;
  assign mem[2982] = 4'h0;
  assign mem[2983] = 4'h3;
  assign mem[2984] = 4'h0;
  assign mem[2985] = 4'h1;
  assign mem[2986] = 4'h0;
  assign mem[2987] = 4'h2;
  assign mem[2988] = 4'h0;
  assign mem[2989] = 4'h1;
  assign mem[2990] = 4'h0;
  assign mem[2991] = 4'h4;
  assign mem[2992] = 4'h0;
  assign mem[2993] = 4'h1;
  assign mem[2994] = 4'h0;
  assign mem[2995] = 4'h2;
  assign mem[2996] = 4'h0;
  assign mem[2997] = 4'h1;
  assign mem[2998] = 4'h0;
  assign mem[2999] = 4'h3;
  assign mem[3000] = 4'h0;
  assign mem[3001] = 4'h1;
  assign mem[3002] = 4'h0;
  assign mem[3003] = 4'h2;
  assign mem[3004] = 4'h0;
  assign mem[3005] = 4'h1;
  assign mem[3006] = 4'h0;
  assign mem[3007] = 4'h6;
  assign mem[3008] = 4'h0;
  assign mem[3009] = 4'h1;
  assign mem[3010] = 4'h0;
  assign mem[3011] = 4'h2;
  assign mem[3012] = 4'h0;
  assign mem[3013] = 4'h1;
  assign mem[3014] = 4'h0;
  assign mem[3015] = 4'h3;
  assign mem[3016] = 4'h0;
  assign mem[3017] = 4'h1;
  assign mem[3018] = 4'h0;
  assign mem[3019] = 4'h2;
  assign mem[3020] = 4'h0;
  assign mem[3021] = 4'h1;
  assign mem[3022] = 4'h0;
  assign mem[3023] = 4'h4;
  assign mem[3024] = 4'h0;
  assign mem[3025] = 4'h1;
  assign mem[3026] = 4'h0;
  assign mem[3027] = 4'h2;
  assign mem[3028] = 4'h0;
  assign mem[3029] = 4'h1;
  assign mem[3030] = 4'h0;
  assign mem[3031] = 4'h3;
  assign mem[3032] = 4'h0;
  assign mem[3033] = 4'h1;
  assign mem[3034] = 4'h0;
  assign mem[3035] = 4'h2;
  assign mem[3036] = 4'h0;
  assign mem[3037] = 4'h1;
  assign mem[3038] = 4'h0;
  assign mem[3039] = 4'h5;
  assign mem[3040] = 4'h0;
  assign mem[3041] = 4'h1;
  assign mem[3042] = 4'h0;
  assign mem[3043] = 4'h2;
  assign mem[3044] = 4'h0;
  assign mem[3045] = 4'h1;
  assign mem[3046] = 4'h0;
  assign mem[3047] = 4'h3;
  assign mem[3048] = 4'h0;
  assign mem[3049] = 4'h1;
  assign mem[3050] = 4'h0;
  assign mem[3051] = 4'h2;
  assign mem[3052] = 4'h0;
  assign mem[3053] = 4'h1;
  assign mem[3054] = 4'h0;
  assign mem[3055] = 4'h4;
  assign mem[3056] = 4'h0;
  assign mem[3057] = 4'h1;
  assign mem[3058] = 4'h0;
  assign mem[3059] = 4'h2;
  assign mem[3060] = 4'h0;
  assign mem[3061] = 4'h1;
  assign mem[3062] = 4'h0;
  assign mem[3063] = 4'h3;
  assign mem[3064] = 4'h0;
  assign mem[3065] = 4'h1;
  assign mem[3066] = 4'h0;
  assign mem[3067] = 4'h2;
  assign mem[3068] = 4'h0;
  assign mem[3069] = 4'h1;
  assign mem[3070] = 4'h0;
  assign mem[3071] = 4'ha;
  assign mem[3072] = 4'h0;
  assign mem[3073] = 4'h1;
  assign mem[3074] = 4'h0;
  assign mem[3075] = 4'h2;
  assign mem[3076] = 4'h0;
  assign mem[3077] = 4'h1;
  assign mem[3078] = 4'h0;
  assign mem[3079] = 4'h3;
  assign mem[3080] = 4'h0;
  assign mem[3081] = 4'h1;
  assign mem[3082] = 4'h0;
  assign mem[3083] = 4'h2;
  assign mem[3084] = 4'h0;
  assign mem[3085] = 4'h1;
  assign mem[3086] = 4'h0;
  assign mem[3087] = 4'h4;
  assign mem[3088] = 4'h0;
  assign mem[3089] = 4'h1;
  assign mem[3090] = 4'h0;
  assign mem[3091] = 4'h2;
  assign mem[3092] = 4'h0;
  assign mem[3093] = 4'h1;
  assign mem[3094] = 4'h0;
  assign mem[3095] = 4'h3;
  assign mem[3096] = 4'h0;
  assign mem[3097] = 4'h1;
  assign mem[3098] = 4'h0;
  assign mem[3099] = 4'h2;
  assign mem[3100] = 4'h0;
  assign mem[3101] = 4'h1;
  assign mem[3102] = 4'h0;
  assign mem[3103] = 4'h5;
  assign mem[3104] = 4'h0;
  assign mem[3105] = 4'h1;
  assign mem[3106] = 4'h0;
  assign mem[3107] = 4'h2;
  assign mem[3108] = 4'h0;
  assign mem[3109] = 4'h1;
  assign mem[3110] = 4'h0;
  assign mem[3111] = 4'h3;
  assign mem[3112] = 4'h0;
  assign mem[3113] = 4'h1;
  assign mem[3114] = 4'h0;
  assign mem[3115] = 4'h2;
  assign mem[3116] = 4'h0;
  assign mem[3117] = 4'h1;
  assign mem[3118] = 4'h0;
  assign mem[3119] = 4'h4;
  assign mem[3120] = 4'h0;
  assign mem[3121] = 4'h1;
  assign mem[3122] = 4'h0;
  assign mem[3123] = 4'h2;
  assign mem[3124] = 4'h0;
  assign mem[3125] = 4'h1;
  assign mem[3126] = 4'h0;
  assign mem[3127] = 4'h3;
  assign mem[3128] = 4'h0;
  assign mem[3129] = 4'h1;
  assign mem[3130] = 4'h0;
  assign mem[3131] = 4'h2;
  assign mem[3132] = 4'h0;
  assign mem[3133] = 4'h1;
  assign mem[3134] = 4'h0;
  assign mem[3135] = 4'h6;
  assign mem[3136] = 4'h0;
  assign mem[3137] = 4'h1;
  assign mem[3138] = 4'h0;
  assign mem[3139] = 4'h2;
  assign mem[3140] = 4'h0;
  assign mem[3141] = 4'h1;
  assign mem[3142] = 4'h0;
  assign mem[3143] = 4'h3;
  assign mem[3144] = 4'h0;
  assign mem[3145] = 4'h1;
  assign mem[3146] = 4'h0;
  assign mem[3147] = 4'h2;
  assign mem[3148] = 4'h0;
  assign mem[3149] = 4'h1;
  assign mem[3150] = 4'h0;
  assign mem[3151] = 4'h4;
  assign mem[3152] = 4'h0;
  assign mem[3153] = 4'h1;
  assign mem[3154] = 4'h0;
  assign mem[3155] = 4'h2;
  assign mem[3156] = 4'h0;
  assign mem[3157] = 4'h1;
  assign mem[3158] = 4'h0;
  assign mem[3159] = 4'h3;
  assign mem[3160] = 4'h0;
  assign mem[3161] = 4'h1;
  assign mem[3162] = 4'h0;
  assign mem[3163] = 4'h2;
  assign mem[3164] = 4'h0;
  assign mem[3165] = 4'h1;
  assign mem[3166] = 4'h0;
  assign mem[3167] = 4'h5;
  assign mem[3168] = 4'h0;
  assign mem[3169] = 4'h1;
  assign mem[3170] = 4'h0;
  assign mem[3171] = 4'h2;
  assign mem[3172] = 4'h0;
  assign mem[3173] = 4'h1;
  assign mem[3174] = 4'h0;
  assign mem[3175] = 4'h3;
  assign mem[3176] = 4'h0;
  assign mem[3177] = 4'h1;
  assign mem[3178] = 4'h0;
  assign mem[3179] = 4'h2;
  assign mem[3180] = 4'h0;
  assign mem[3181] = 4'h1;
  assign mem[3182] = 4'h0;
  assign mem[3183] = 4'h4;
  assign mem[3184] = 4'h0;
  assign mem[3185] = 4'h1;
  assign mem[3186] = 4'h0;
  assign mem[3187] = 4'h2;
  assign mem[3188] = 4'h0;
  assign mem[3189] = 4'h1;
  assign mem[3190] = 4'h0;
  assign mem[3191] = 4'h3;
  assign mem[3192] = 4'h0;
  assign mem[3193] = 4'h1;
  assign mem[3194] = 4'h0;
  assign mem[3195] = 4'h2;
  assign mem[3196] = 4'h0;
  assign mem[3197] = 4'h1;
  assign mem[3198] = 4'h0;
  assign mem[3199] = 4'h7;
  assign mem[3200] = 4'h0;
  assign mem[3201] = 4'h1;
  assign mem[3202] = 4'h0;
  assign mem[3203] = 4'h2;
  assign mem[3204] = 4'h0;
  assign mem[3205] = 4'h1;
  assign mem[3206] = 4'h0;
  assign mem[3207] = 4'h3;
  assign mem[3208] = 4'h0;
  assign mem[3209] = 4'h1;
  assign mem[3210] = 4'h0;
  assign mem[3211] = 4'h2;
  assign mem[3212] = 4'h0;
  assign mem[3213] = 4'h1;
  assign mem[3214] = 4'h0;
  assign mem[3215] = 4'h4;
  assign mem[3216] = 4'h0;
  assign mem[3217] = 4'h1;
  assign mem[3218] = 4'h0;
  assign mem[3219] = 4'h2;
  assign mem[3220] = 4'h0;
  assign mem[3221] = 4'h1;
  assign mem[3222] = 4'h0;
  assign mem[3223] = 4'h3;
  assign mem[3224] = 4'h0;
  assign mem[3225] = 4'h1;
  assign mem[3226] = 4'h0;
  assign mem[3227] = 4'h2;
  assign mem[3228] = 4'h0;
  assign mem[3229] = 4'h1;
  assign mem[3230] = 4'h0;
  assign mem[3231] = 4'h5;
  assign mem[3232] = 4'h0;
  assign mem[3233] = 4'h1;
  assign mem[3234] = 4'h0;
  assign mem[3235] = 4'h2;
  assign mem[3236] = 4'h0;
  assign mem[3237] = 4'h1;
  assign mem[3238] = 4'h0;
  assign mem[3239] = 4'h3;
  assign mem[3240] = 4'h0;
  assign mem[3241] = 4'h1;
  assign mem[3242] = 4'h0;
  assign mem[3243] = 4'h2;
  assign mem[3244] = 4'h0;
  assign mem[3245] = 4'h1;
  assign mem[3246] = 4'h0;
  assign mem[3247] = 4'h4;
  assign mem[3248] = 4'h0;
  assign mem[3249] = 4'h1;
  assign mem[3250] = 4'h0;
  assign mem[3251] = 4'h2;
  assign mem[3252] = 4'h0;
  assign mem[3253] = 4'h1;
  assign mem[3254] = 4'h0;
  assign mem[3255] = 4'h3;
  assign mem[3256] = 4'h0;
  assign mem[3257] = 4'h1;
  assign mem[3258] = 4'h0;
  assign mem[3259] = 4'h2;
  assign mem[3260] = 4'h0;
  assign mem[3261] = 4'h1;
  assign mem[3262] = 4'h0;
  assign mem[3263] = 4'h6;
  assign mem[3264] = 4'h0;
  assign mem[3265] = 4'h1;
  assign mem[3266] = 4'h0;
  assign mem[3267] = 4'h2;
  assign mem[3268] = 4'h0;
  assign mem[3269] = 4'h1;
  assign mem[3270] = 4'h0;
  assign mem[3271] = 4'h3;
  assign mem[3272] = 4'h0;
  assign mem[3273] = 4'h1;
  assign mem[3274] = 4'h0;
  assign mem[3275] = 4'h2;
  assign mem[3276] = 4'h0;
  assign mem[3277] = 4'h1;
  assign mem[3278] = 4'h0;
  assign mem[3279] = 4'h4;
  assign mem[3280] = 4'h0;
  assign mem[3281] = 4'h1;
  assign mem[3282] = 4'h0;
  assign mem[3283] = 4'h2;
  assign mem[3284] = 4'h0;
  assign mem[3285] = 4'h1;
  assign mem[3286] = 4'h0;
  assign mem[3287] = 4'h3;
  assign mem[3288] = 4'h0;
  assign mem[3289] = 4'h1;
  assign mem[3290] = 4'h0;
  assign mem[3291] = 4'h2;
  assign mem[3292] = 4'h0;
  assign mem[3293] = 4'h1;
  assign mem[3294] = 4'h0;
  assign mem[3295] = 4'h5;
  assign mem[3296] = 4'h0;
  assign mem[3297] = 4'h1;
  assign mem[3298] = 4'h0;
  assign mem[3299] = 4'h2;
  assign mem[3300] = 4'h0;
  assign mem[3301] = 4'h1;
  assign mem[3302] = 4'h0;
  assign mem[3303] = 4'h3;
  assign mem[3304] = 4'h0;
  assign mem[3305] = 4'h1;
  assign mem[3306] = 4'h0;
  assign mem[3307] = 4'h2;
  assign mem[3308] = 4'h0;
  assign mem[3309] = 4'h1;
  assign mem[3310] = 4'h0;
  assign mem[3311] = 4'h4;
  assign mem[3312] = 4'h0;
  assign mem[3313] = 4'h1;
  assign mem[3314] = 4'h0;
  assign mem[3315] = 4'h2;
  assign mem[3316] = 4'h0;
  assign mem[3317] = 4'h1;
  assign mem[3318] = 4'h0;
  assign mem[3319] = 4'h3;
  assign mem[3320] = 4'h0;
  assign mem[3321] = 4'h1;
  assign mem[3322] = 4'h0;
  assign mem[3323] = 4'h2;
  assign mem[3324] = 4'h0;
  assign mem[3325] = 4'h1;
  assign mem[3326] = 4'h0;
  assign mem[3327] = 4'h8;
  assign mem[3328] = 4'h0;
  assign mem[3329] = 4'h1;
  assign mem[3330] = 4'h0;
  assign mem[3331] = 4'h2;
  assign mem[3332] = 4'h0;
  assign mem[3333] = 4'h1;
  assign mem[3334] = 4'h0;
  assign mem[3335] = 4'h3;
  assign mem[3336] = 4'h0;
  assign mem[3337] = 4'h1;
  assign mem[3338] = 4'h0;
  assign mem[3339] = 4'h2;
  assign mem[3340] = 4'h0;
  assign mem[3341] = 4'h1;
  assign mem[3342] = 4'h0;
  assign mem[3343] = 4'h4;
  assign mem[3344] = 4'h0;
  assign mem[3345] = 4'h1;
  assign mem[3346] = 4'h0;
  assign mem[3347] = 4'h2;
  assign mem[3348] = 4'h0;
  assign mem[3349] = 4'h1;
  assign mem[3350] = 4'h0;
  assign mem[3351] = 4'h3;
  assign mem[3352] = 4'h0;
  assign mem[3353] = 4'h1;
  assign mem[3354] = 4'h0;
  assign mem[3355] = 4'h2;
  assign mem[3356] = 4'h0;
  assign mem[3357] = 4'h1;
  assign mem[3358] = 4'h0;
  assign mem[3359] = 4'h5;
  assign mem[3360] = 4'h0;
  assign mem[3361] = 4'h1;
  assign mem[3362] = 4'h0;
  assign mem[3363] = 4'h2;
  assign mem[3364] = 4'h0;
  assign mem[3365] = 4'h1;
  assign mem[3366] = 4'h0;
  assign mem[3367] = 4'h3;
  assign mem[3368] = 4'h0;
  assign mem[3369] = 4'h1;
  assign mem[3370] = 4'h0;
  assign mem[3371] = 4'h2;
  assign mem[3372] = 4'h0;
  assign mem[3373] = 4'h1;
  assign mem[3374] = 4'h0;
  assign mem[3375] = 4'h4;
  assign mem[3376] = 4'h0;
  assign mem[3377] = 4'h1;
  assign mem[3378] = 4'h0;
  assign mem[3379] = 4'h2;
  assign mem[3380] = 4'h0;
  assign mem[3381] = 4'h1;
  assign mem[3382] = 4'h0;
  assign mem[3383] = 4'h3;
  assign mem[3384] = 4'h0;
  assign mem[3385] = 4'h1;
  assign mem[3386] = 4'h0;
  assign mem[3387] = 4'h2;
  assign mem[3388] = 4'h0;
  assign mem[3389] = 4'h1;
  assign mem[3390] = 4'h0;
  assign mem[3391] = 4'h6;
  assign mem[3392] = 4'h0;
  assign mem[3393] = 4'h1;
  assign mem[3394] = 4'h0;
  assign mem[3395] = 4'h2;
  assign mem[3396] = 4'h0;
  assign mem[3397] = 4'h1;
  assign mem[3398] = 4'h0;
  assign mem[3399] = 4'h3;
  assign mem[3400] = 4'h0;
  assign mem[3401] = 4'h1;
  assign mem[3402] = 4'h0;
  assign mem[3403] = 4'h2;
  assign mem[3404] = 4'h0;
  assign mem[3405] = 4'h1;
  assign mem[3406] = 4'h0;
  assign mem[3407] = 4'h4;
  assign mem[3408] = 4'h0;
  assign mem[3409] = 4'h1;
  assign mem[3410] = 4'h0;
  assign mem[3411] = 4'h2;
  assign mem[3412] = 4'h0;
  assign mem[3413] = 4'h1;
  assign mem[3414] = 4'h0;
  assign mem[3415] = 4'h3;
  assign mem[3416] = 4'h0;
  assign mem[3417] = 4'h1;
  assign mem[3418] = 4'h0;
  assign mem[3419] = 4'h2;
  assign mem[3420] = 4'h0;
  assign mem[3421] = 4'h1;
  assign mem[3422] = 4'h0;
  assign mem[3423] = 4'h5;
  assign mem[3424] = 4'h0;
  assign mem[3425] = 4'h1;
  assign mem[3426] = 4'h0;
  assign mem[3427] = 4'h2;
  assign mem[3428] = 4'h0;
  assign mem[3429] = 4'h1;
  assign mem[3430] = 4'h0;
  assign mem[3431] = 4'h3;
  assign mem[3432] = 4'h0;
  assign mem[3433] = 4'h1;
  assign mem[3434] = 4'h0;
  assign mem[3435] = 4'h2;
  assign mem[3436] = 4'h0;
  assign mem[3437] = 4'h1;
  assign mem[3438] = 4'h0;
  assign mem[3439] = 4'h4;
  assign mem[3440] = 4'h0;
  assign mem[3441] = 4'h1;
  assign mem[3442] = 4'h0;
  assign mem[3443] = 4'h2;
  assign mem[3444] = 4'h0;
  assign mem[3445] = 4'h1;
  assign mem[3446] = 4'h0;
  assign mem[3447] = 4'h3;
  assign mem[3448] = 4'h0;
  assign mem[3449] = 4'h1;
  assign mem[3450] = 4'h0;
  assign mem[3451] = 4'h2;
  assign mem[3452] = 4'h0;
  assign mem[3453] = 4'h1;
  assign mem[3454] = 4'h0;
  assign mem[3455] = 4'h7;
  assign mem[3456] = 4'h0;
  assign mem[3457] = 4'h1;
  assign mem[3458] = 4'h0;
  assign mem[3459] = 4'h2;
  assign mem[3460] = 4'h0;
  assign mem[3461] = 4'h1;
  assign mem[3462] = 4'h0;
  assign mem[3463] = 4'h3;
  assign mem[3464] = 4'h0;
  assign mem[3465] = 4'h1;
  assign mem[3466] = 4'h0;
  assign mem[3467] = 4'h2;
  assign mem[3468] = 4'h0;
  assign mem[3469] = 4'h1;
  assign mem[3470] = 4'h0;
  assign mem[3471] = 4'h4;
  assign mem[3472] = 4'h0;
  assign mem[3473] = 4'h1;
  assign mem[3474] = 4'h0;
  assign mem[3475] = 4'h2;
  assign mem[3476] = 4'h0;
  assign mem[3477] = 4'h1;
  assign mem[3478] = 4'h0;
  assign mem[3479] = 4'h3;
  assign mem[3480] = 4'h0;
  assign mem[3481] = 4'h1;
  assign mem[3482] = 4'h0;
  assign mem[3483] = 4'h2;
  assign mem[3484] = 4'h0;
  assign mem[3485] = 4'h1;
  assign mem[3486] = 4'h0;
  assign mem[3487] = 4'h5;
  assign mem[3488] = 4'h0;
  assign mem[3489] = 4'h1;
  assign mem[3490] = 4'h0;
  assign mem[3491] = 4'h2;
  assign mem[3492] = 4'h0;
  assign mem[3493] = 4'h1;
  assign mem[3494] = 4'h0;
  assign mem[3495] = 4'h3;
  assign mem[3496] = 4'h0;
  assign mem[3497] = 4'h1;
  assign mem[3498] = 4'h0;
  assign mem[3499] = 4'h2;
  assign mem[3500] = 4'h0;
  assign mem[3501] = 4'h1;
  assign mem[3502] = 4'h0;
  assign mem[3503] = 4'h4;
  assign mem[3504] = 4'h0;
  assign mem[3505] = 4'h1;
  assign mem[3506] = 4'h0;
  assign mem[3507] = 4'h2;
  assign mem[3508] = 4'h0;
  assign mem[3509] = 4'h1;
  assign mem[3510] = 4'h0;
  assign mem[3511] = 4'h3;
  assign mem[3512] = 4'h0;
  assign mem[3513] = 4'h1;
  assign mem[3514] = 4'h0;
  assign mem[3515] = 4'h2;
  assign mem[3516] = 4'h0;
  assign mem[3517] = 4'h1;
  assign mem[3518] = 4'h0;
  assign mem[3519] = 4'h6;
  assign mem[3520] = 4'h0;
  assign mem[3521] = 4'h1;
  assign mem[3522] = 4'h0;
  assign mem[3523] = 4'h2;
  assign mem[3524] = 4'h0;
  assign mem[3525] = 4'h1;
  assign mem[3526] = 4'h0;
  assign mem[3527] = 4'h3;
  assign mem[3528] = 4'h0;
  assign mem[3529] = 4'h1;
  assign mem[3530] = 4'h0;
  assign mem[3531] = 4'h2;
  assign mem[3532] = 4'h0;
  assign mem[3533] = 4'h1;
  assign mem[3534] = 4'h0;
  assign mem[3535] = 4'h4;
  assign mem[3536] = 4'h0;
  assign mem[3537] = 4'h1;
  assign mem[3538] = 4'h0;
  assign mem[3539] = 4'h2;
  assign mem[3540] = 4'h0;
  assign mem[3541] = 4'h1;
  assign mem[3542] = 4'h0;
  assign mem[3543] = 4'h3;
  assign mem[3544] = 4'h0;
  assign mem[3545] = 4'h1;
  assign mem[3546] = 4'h0;
  assign mem[3547] = 4'h2;
  assign mem[3548] = 4'h0;
  assign mem[3549] = 4'h1;
  assign mem[3550] = 4'h0;
  assign mem[3551] = 4'h5;
  assign mem[3552] = 4'h0;
  assign mem[3553] = 4'h1;
  assign mem[3554] = 4'h0;
  assign mem[3555] = 4'h2;
  assign mem[3556] = 4'h0;
  assign mem[3557] = 4'h1;
  assign mem[3558] = 4'h0;
  assign mem[3559] = 4'h3;
  assign mem[3560] = 4'h0;
  assign mem[3561] = 4'h1;
  assign mem[3562] = 4'h0;
  assign mem[3563] = 4'h2;
  assign mem[3564] = 4'h0;
  assign mem[3565] = 4'h1;
  assign mem[3566] = 4'h0;
  assign mem[3567] = 4'h4;
  assign mem[3568] = 4'h0;
  assign mem[3569] = 4'h1;
  assign mem[3570] = 4'h0;
  assign mem[3571] = 4'h2;
  assign mem[3572] = 4'h0;
  assign mem[3573] = 4'h1;
  assign mem[3574] = 4'h0;
  assign mem[3575] = 4'h3;
  assign mem[3576] = 4'h0;
  assign mem[3577] = 4'h1;
  assign mem[3578] = 4'h0;
  assign mem[3579] = 4'h2;
  assign mem[3580] = 4'h0;
  assign mem[3581] = 4'h1;
  assign mem[3582] = 4'h0;
  assign mem[3583] = 4'h9;
  assign mem[3584] = 4'h0;
  assign mem[3585] = 4'h1;
  assign mem[3586] = 4'h0;
  assign mem[3587] = 4'h2;
  assign mem[3588] = 4'h0;
  assign mem[3589] = 4'h1;
  assign mem[3590] = 4'h0;
  assign mem[3591] = 4'h3;
  assign mem[3592] = 4'h0;
  assign mem[3593] = 4'h1;
  assign mem[3594] = 4'h0;
  assign mem[3595] = 4'h2;
  assign mem[3596] = 4'h0;
  assign mem[3597] = 4'h1;
  assign mem[3598] = 4'h0;
  assign mem[3599] = 4'h4;
  assign mem[3600] = 4'h0;
  assign mem[3601] = 4'h1;
  assign mem[3602] = 4'h0;
  assign mem[3603] = 4'h2;
  assign mem[3604] = 4'h0;
  assign mem[3605] = 4'h1;
  assign mem[3606] = 4'h0;
  assign mem[3607] = 4'h3;
  assign mem[3608] = 4'h0;
  assign mem[3609] = 4'h1;
  assign mem[3610] = 4'h0;
  assign mem[3611] = 4'h2;
  assign mem[3612] = 4'h0;
  assign mem[3613] = 4'h1;
  assign mem[3614] = 4'h0;
  assign mem[3615] = 4'h5;
  assign mem[3616] = 4'h0;
  assign mem[3617] = 4'h1;
  assign mem[3618] = 4'h0;
  assign mem[3619] = 4'h2;
  assign mem[3620] = 4'h0;
  assign mem[3621] = 4'h1;
  assign mem[3622] = 4'h0;
  assign mem[3623] = 4'h3;
  assign mem[3624] = 4'h0;
  assign mem[3625] = 4'h1;
  assign mem[3626] = 4'h0;
  assign mem[3627] = 4'h2;
  assign mem[3628] = 4'h0;
  assign mem[3629] = 4'h1;
  assign mem[3630] = 4'h0;
  assign mem[3631] = 4'h4;
  assign mem[3632] = 4'h0;
  assign mem[3633] = 4'h1;
  assign mem[3634] = 4'h0;
  assign mem[3635] = 4'h2;
  assign mem[3636] = 4'h0;
  assign mem[3637] = 4'h1;
  assign mem[3638] = 4'h0;
  assign mem[3639] = 4'h3;
  assign mem[3640] = 4'h0;
  assign mem[3641] = 4'h1;
  assign mem[3642] = 4'h0;
  assign mem[3643] = 4'h2;
  assign mem[3644] = 4'h0;
  assign mem[3645] = 4'h1;
  assign mem[3646] = 4'h0;
  assign mem[3647] = 4'h6;
  assign mem[3648] = 4'h0;
  assign mem[3649] = 4'h1;
  assign mem[3650] = 4'h0;
  assign mem[3651] = 4'h2;
  assign mem[3652] = 4'h0;
  assign mem[3653] = 4'h1;
  assign mem[3654] = 4'h0;
  assign mem[3655] = 4'h3;
  assign mem[3656] = 4'h0;
  assign mem[3657] = 4'h1;
  assign mem[3658] = 4'h0;
  assign mem[3659] = 4'h2;
  assign mem[3660] = 4'h0;
  assign mem[3661] = 4'h1;
  assign mem[3662] = 4'h0;
  assign mem[3663] = 4'h4;
  assign mem[3664] = 4'h0;
  assign mem[3665] = 4'h1;
  assign mem[3666] = 4'h0;
  assign mem[3667] = 4'h2;
  assign mem[3668] = 4'h0;
  assign mem[3669] = 4'h1;
  assign mem[3670] = 4'h0;
  assign mem[3671] = 4'h3;
  assign mem[3672] = 4'h0;
  assign mem[3673] = 4'h1;
  assign mem[3674] = 4'h0;
  assign mem[3675] = 4'h2;
  assign mem[3676] = 4'h0;
  assign mem[3677] = 4'h1;
  assign mem[3678] = 4'h0;
  assign mem[3679] = 4'h5;
  assign mem[3680] = 4'h0;
  assign mem[3681] = 4'h1;
  assign mem[3682] = 4'h0;
  assign mem[3683] = 4'h2;
  assign mem[3684] = 4'h0;
  assign mem[3685] = 4'h1;
  assign mem[3686] = 4'h0;
  assign mem[3687] = 4'h3;
  assign mem[3688] = 4'h0;
  assign mem[3689] = 4'h1;
  assign mem[3690] = 4'h0;
  assign mem[3691] = 4'h2;
  assign mem[3692] = 4'h0;
  assign mem[3693] = 4'h1;
  assign mem[3694] = 4'h0;
  assign mem[3695] = 4'h4;
  assign mem[3696] = 4'h0;
  assign mem[3697] = 4'h1;
  assign mem[3698] = 4'h0;
  assign mem[3699] = 4'h2;
  assign mem[3700] = 4'h0;
  assign mem[3701] = 4'h1;
  assign mem[3702] = 4'h0;
  assign mem[3703] = 4'h3;
  assign mem[3704] = 4'h0;
  assign mem[3705] = 4'h1;
  assign mem[3706] = 4'h0;
  assign mem[3707] = 4'h2;
  assign mem[3708] = 4'h0;
  assign mem[3709] = 4'h1;
  assign mem[3710] = 4'h0;
  assign mem[3711] = 4'h7;
  assign mem[3712] = 4'h0;
  assign mem[3713] = 4'h1;
  assign mem[3714] = 4'h0;
  assign mem[3715] = 4'h2;
  assign mem[3716] = 4'h0;
  assign mem[3717] = 4'h1;
  assign mem[3718] = 4'h0;
  assign mem[3719] = 4'h3;
  assign mem[3720] = 4'h0;
  assign mem[3721] = 4'h1;
  assign mem[3722] = 4'h0;
  assign mem[3723] = 4'h2;
  assign mem[3724] = 4'h0;
  assign mem[3725] = 4'h1;
  assign mem[3726] = 4'h0;
  assign mem[3727] = 4'h4;
  assign mem[3728] = 4'h0;
  assign mem[3729] = 4'h1;
  assign mem[3730] = 4'h0;
  assign mem[3731] = 4'h2;
  assign mem[3732] = 4'h0;
  assign mem[3733] = 4'h1;
  assign mem[3734] = 4'h0;
  assign mem[3735] = 4'h3;
  assign mem[3736] = 4'h0;
  assign mem[3737] = 4'h1;
  assign mem[3738] = 4'h0;
  assign mem[3739] = 4'h2;
  assign mem[3740] = 4'h0;
  assign mem[3741] = 4'h1;
  assign mem[3742] = 4'h0;
  assign mem[3743] = 4'h5;
  assign mem[3744] = 4'h0;
  assign mem[3745] = 4'h1;
  assign mem[3746] = 4'h0;
  assign mem[3747] = 4'h2;
  assign mem[3748] = 4'h0;
  assign mem[3749] = 4'h1;
  assign mem[3750] = 4'h0;
  assign mem[3751] = 4'h3;
  assign mem[3752] = 4'h0;
  assign mem[3753] = 4'h1;
  assign mem[3754] = 4'h0;
  assign mem[3755] = 4'h2;
  assign mem[3756] = 4'h0;
  assign mem[3757] = 4'h1;
  assign mem[3758] = 4'h0;
  assign mem[3759] = 4'h4;
  assign mem[3760] = 4'h0;
  assign mem[3761] = 4'h1;
  assign mem[3762] = 4'h0;
  assign mem[3763] = 4'h2;
  assign mem[3764] = 4'h0;
  assign mem[3765] = 4'h1;
  assign mem[3766] = 4'h0;
  assign mem[3767] = 4'h3;
  assign mem[3768] = 4'h0;
  assign mem[3769] = 4'h1;
  assign mem[3770] = 4'h0;
  assign mem[3771] = 4'h2;
  assign mem[3772] = 4'h0;
  assign mem[3773] = 4'h1;
  assign mem[3774] = 4'h0;
  assign mem[3775] = 4'h6;
  assign mem[3776] = 4'h0;
  assign mem[3777] = 4'h1;
  assign mem[3778] = 4'h0;
  assign mem[3779] = 4'h2;
  assign mem[3780] = 4'h0;
  assign mem[3781] = 4'h1;
  assign mem[3782] = 4'h0;
  assign mem[3783] = 4'h3;
  assign mem[3784] = 4'h0;
  assign mem[3785] = 4'h1;
  assign mem[3786] = 4'h0;
  assign mem[3787] = 4'h2;
  assign mem[3788] = 4'h0;
  assign mem[3789] = 4'h1;
  assign mem[3790] = 4'h0;
  assign mem[3791] = 4'h4;
  assign mem[3792] = 4'h0;
  assign mem[3793] = 4'h1;
  assign mem[3794] = 4'h0;
  assign mem[3795] = 4'h2;
  assign mem[3796] = 4'h0;
  assign mem[3797] = 4'h1;
  assign mem[3798] = 4'h0;
  assign mem[3799] = 4'h3;
  assign mem[3800] = 4'h0;
  assign mem[3801] = 4'h1;
  assign mem[3802] = 4'h0;
  assign mem[3803] = 4'h2;
  assign mem[3804] = 4'h0;
  assign mem[3805] = 4'h1;
  assign mem[3806] = 4'h0;
  assign mem[3807] = 4'h5;
  assign mem[3808] = 4'h0;
  assign mem[3809] = 4'h1;
  assign mem[3810] = 4'h0;
  assign mem[3811] = 4'h2;
  assign mem[3812] = 4'h0;
  assign mem[3813] = 4'h1;
  assign mem[3814] = 4'h0;
  assign mem[3815] = 4'h3;
  assign mem[3816] = 4'h0;
  assign mem[3817] = 4'h1;
  assign mem[3818] = 4'h0;
  assign mem[3819] = 4'h2;
  assign mem[3820] = 4'h0;
  assign mem[3821] = 4'h1;
  assign mem[3822] = 4'h0;
  assign mem[3823] = 4'h4;
  assign mem[3824] = 4'h0;
  assign mem[3825] = 4'h1;
  assign mem[3826] = 4'h0;
  assign mem[3827] = 4'h2;
  assign mem[3828] = 4'h0;
  assign mem[3829] = 4'h1;
  assign mem[3830] = 4'h0;
  assign mem[3831] = 4'h3;
  assign mem[3832] = 4'h0;
  assign mem[3833] = 4'h1;
  assign mem[3834] = 4'h0;
  assign mem[3835] = 4'h2;
  assign mem[3836] = 4'h0;
  assign mem[3837] = 4'h1;
  assign mem[3838] = 4'h0;
  assign mem[3839] = 4'h8;
  assign mem[3840] = 4'h0;
  assign mem[3841] = 4'h1;
  assign mem[3842] = 4'h0;
  assign mem[3843] = 4'h2;
  assign mem[3844] = 4'h0;
  assign mem[3845] = 4'h1;
  assign mem[3846] = 4'h0;
  assign mem[3847] = 4'h3;
  assign mem[3848] = 4'h0;
  assign mem[3849] = 4'h1;
  assign mem[3850] = 4'h0;
  assign mem[3851] = 4'h2;
  assign mem[3852] = 4'h0;
  assign mem[3853] = 4'h1;
  assign mem[3854] = 4'h0;
  assign mem[3855] = 4'h4;
  assign mem[3856] = 4'h0;
  assign mem[3857] = 4'h1;
  assign mem[3858] = 4'h0;
  assign mem[3859] = 4'h2;
  assign mem[3860] = 4'h0;
  assign mem[3861] = 4'h1;
  assign mem[3862] = 4'h0;
  assign mem[3863] = 4'h3;
  assign mem[3864] = 4'h0;
  assign mem[3865] = 4'h1;
  assign mem[3866] = 4'h0;
  assign mem[3867] = 4'h2;
  assign mem[3868] = 4'h0;
  assign mem[3869] = 4'h1;
  assign mem[3870] = 4'h0;
  assign mem[3871] = 4'h5;
  assign mem[3872] = 4'h0;
  assign mem[3873] = 4'h1;
  assign mem[3874] = 4'h0;
  assign mem[3875] = 4'h2;
  assign mem[3876] = 4'h0;
  assign mem[3877] = 4'h1;
  assign mem[3878] = 4'h0;
  assign mem[3879] = 4'h3;
  assign mem[3880] = 4'h0;
  assign mem[3881] = 4'h1;
  assign mem[3882] = 4'h0;
  assign mem[3883] = 4'h2;
  assign mem[3884] = 4'h0;
  assign mem[3885] = 4'h1;
  assign mem[3886] = 4'h0;
  assign mem[3887] = 4'h4;
  assign mem[3888] = 4'h0;
  assign mem[3889] = 4'h1;
  assign mem[3890] = 4'h0;
  assign mem[3891] = 4'h2;
  assign mem[3892] = 4'h0;
  assign mem[3893] = 4'h1;
  assign mem[3894] = 4'h0;
  assign mem[3895] = 4'h3;
  assign mem[3896] = 4'h0;
  assign mem[3897] = 4'h1;
  assign mem[3898] = 4'h0;
  assign mem[3899] = 4'h2;
  assign mem[3900] = 4'h0;
  assign mem[3901] = 4'h1;
  assign mem[3902] = 4'h0;
  assign mem[3903] = 4'h6;
  assign mem[3904] = 4'h0;
  assign mem[3905] = 4'h1;
  assign mem[3906] = 4'h0;
  assign mem[3907] = 4'h2;
  assign mem[3908] = 4'h0;
  assign mem[3909] = 4'h1;
  assign mem[3910] = 4'h0;
  assign mem[3911] = 4'h3;
  assign mem[3912] = 4'h0;
  assign mem[3913] = 4'h1;
  assign mem[3914] = 4'h0;
  assign mem[3915] = 4'h2;
  assign mem[3916] = 4'h0;
  assign mem[3917] = 4'h1;
  assign mem[3918] = 4'h0;
  assign mem[3919] = 4'h4;
  assign mem[3920] = 4'h0;
  assign mem[3921] = 4'h1;
  assign mem[3922] = 4'h0;
  assign mem[3923] = 4'h2;
  assign mem[3924] = 4'h0;
  assign mem[3925] = 4'h1;
  assign mem[3926] = 4'h0;
  assign mem[3927] = 4'h3;
  assign mem[3928] = 4'h0;
  assign mem[3929] = 4'h1;
  assign mem[3930] = 4'h0;
  assign mem[3931] = 4'h2;
  assign mem[3932] = 4'h0;
  assign mem[3933] = 4'h1;
  assign mem[3934] = 4'h0;
  assign mem[3935] = 4'h5;
  assign mem[3936] = 4'h0;
  assign mem[3937] = 4'h1;
  assign mem[3938] = 4'h0;
  assign mem[3939] = 4'h2;
  assign mem[3940] = 4'h0;
  assign mem[3941] = 4'h1;
  assign mem[3942] = 4'h0;
  assign mem[3943] = 4'h3;
  assign mem[3944] = 4'h0;
  assign mem[3945] = 4'h1;
  assign mem[3946] = 4'h0;
  assign mem[3947] = 4'h2;
  assign mem[3948] = 4'h0;
  assign mem[3949] = 4'h1;
  assign mem[3950] = 4'h0;
  assign mem[3951] = 4'h4;
  assign mem[3952] = 4'h0;
  assign mem[3953] = 4'h1;
  assign mem[3954] = 4'h0;
  assign mem[3955] = 4'h2;
  assign mem[3956] = 4'h0;
  assign mem[3957] = 4'h1;
  assign mem[3958] = 4'h0;
  assign mem[3959] = 4'h3;
  assign mem[3960] = 4'h0;
  assign mem[3961] = 4'h1;
  assign mem[3962] = 4'h0;
  assign mem[3963] = 4'h2;
  assign mem[3964] = 4'h0;
  assign mem[3965] = 4'h1;
  assign mem[3966] = 4'h0;
  assign mem[3967] = 4'h7;
  assign mem[3968] = 4'h0;
  assign mem[3969] = 4'h1;
  assign mem[3970] = 4'h0;
  assign mem[3971] = 4'h2;
  assign mem[3972] = 4'h0;
  assign mem[3973] = 4'h1;
  assign mem[3974] = 4'h0;
  assign mem[3975] = 4'h3;
  assign mem[3976] = 4'h0;
  assign mem[3977] = 4'h1;
  assign mem[3978] = 4'h0;
  assign mem[3979] = 4'h2;
  assign mem[3980] = 4'h0;
  assign mem[3981] = 4'h1;
  assign mem[3982] = 4'h0;
  assign mem[3983] = 4'h4;
  assign mem[3984] = 4'h0;
  assign mem[3985] = 4'h1;
  assign mem[3986] = 4'h0;
  assign mem[3987] = 4'h2;
  assign mem[3988] = 4'h0;
  assign mem[3989] = 4'h1;
  assign mem[3990] = 4'h0;
  assign mem[3991] = 4'h3;
  assign mem[3992] = 4'h0;
  assign mem[3993] = 4'h1;
  assign mem[3994] = 4'h0;
  assign mem[3995] = 4'h2;
  assign mem[3996] = 4'h0;
  assign mem[3997] = 4'h1;
  assign mem[3998] = 4'h0;
  assign mem[3999] = 4'h5;
  assign mem[4000] = 4'h0;
  assign mem[4001] = 4'h1;
  assign mem[4002] = 4'h0;
  assign mem[4003] = 4'h2;
  assign mem[4004] = 4'h0;
  assign mem[4005] = 4'h1;
  assign mem[4006] = 4'h0;
  assign mem[4007] = 4'h3;
  assign mem[4008] = 4'h0;
  assign mem[4009] = 4'h1;
  assign mem[4010] = 4'h0;
  assign mem[4011] = 4'h2;
  assign mem[4012] = 4'h0;
  assign mem[4013] = 4'h1;
  assign mem[4014] = 4'h0;
  assign mem[4015] = 4'h4;
  assign mem[4016] = 4'h0;
  assign mem[4017] = 4'h1;
  assign mem[4018] = 4'h0;
  assign mem[4019] = 4'h2;
  assign mem[4020] = 4'h0;
  assign mem[4021] = 4'h1;
  assign mem[4022] = 4'h0;
  assign mem[4023] = 4'h3;
  assign mem[4024] = 4'h0;
  assign mem[4025] = 4'h1;
  assign mem[4026] = 4'h0;
  assign mem[4027] = 4'h2;
  assign mem[4028] = 4'h0;
  assign mem[4029] = 4'h1;
  assign mem[4030] = 4'h0;
  assign mem[4031] = 4'h6;
  assign mem[4032] = 4'h0;
  assign mem[4033] = 4'h1;
  assign mem[4034] = 4'h0;
  assign mem[4035] = 4'h2;
  assign mem[4036] = 4'h0;
  assign mem[4037] = 4'h1;
  assign mem[4038] = 4'h0;
  assign mem[4039] = 4'h3;
  assign mem[4040] = 4'h0;
  assign mem[4041] = 4'h1;
  assign mem[4042] = 4'h0;
  assign mem[4043] = 4'h2;
  assign mem[4044] = 4'h0;
  assign mem[4045] = 4'h1;
  assign mem[4046] = 4'h0;
  assign mem[4047] = 4'h4;
  assign mem[4048] = 4'h0;
  assign mem[4049] = 4'h1;
  assign mem[4050] = 4'h0;
  assign mem[4051] = 4'h2;
  assign mem[4052] = 4'h0;
  assign mem[4053] = 4'h1;
  assign mem[4054] = 4'h0;
  assign mem[4055] = 4'h3;
  assign mem[4056] = 4'h0;
  assign mem[4057] = 4'h1;
  assign mem[4058] = 4'h0;
  assign mem[4059] = 4'h2;
  assign mem[4060] = 4'h0;
  assign mem[4061] = 4'h1;
  assign mem[4062] = 4'h0;
  assign mem[4063] = 4'h5;
  assign mem[4064] = 4'h0;
  assign mem[4065] = 4'h1;
  assign mem[4066] = 4'h0;
  assign mem[4067] = 4'h2;
  assign mem[4068] = 4'h0;
  assign mem[4069] = 4'h1;
  assign mem[4070] = 4'h0;
  assign mem[4071] = 4'h3;
  assign mem[4072] = 4'h0;
  assign mem[4073] = 4'h1;
  assign mem[4074] = 4'h0;
  assign mem[4075] = 4'h2;
  assign mem[4076] = 4'h0;
  assign mem[4077] = 4'h1;
  assign mem[4078] = 4'h0;
  assign mem[4079] = 4'h4;
  assign mem[4080] = 4'h0;
  assign mem[4081] = 4'h1;
  assign mem[4082] = 4'h0;
  assign mem[4083] = 4'h2;
  assign mem[4084] = 4'h0;
  assign mem[4085] = 4'h1;
  assign mem[4086] = 4'h0;
  assign mem[4087] = 4'h3;
  assign mem[4088] = 4'h0;
  assign mem[4089] = 4'h1;
  assign mem[4090] = 4'h0;
  assign mem[4091] = 4'h2;
  assign mem[4092] = 4'h0;
  assign mem[4093] = 4'h1;
  assign mem[4094] = 4'h0;
  assign mem[4095] = 4'h0; 
  
  //----
  generate 
  if (RD_TYPE==0)
  begin:U_type0
    reg [$clog2(D)-1:0]addr_d1;

    always @(posedge clk)
    begin
      if((!we) & ce)
        addr_d1 <= addr;
    end

    assign rdata = mem[addr_d1];
  end
  else 
  begin:U_type1

    reg [W-1:0]rdata_int;
    always @(posedge clk)
    begin
      if((!we) & ce)
        rdata_int <= mem[addr];
    end

    assign rdata = rdata_int;
  end
  endgenerate
endmodule
