//////////////////////////////////////////////////////////////////////////////////
// Description   : pdec_reg_dyn_bd regfile cfg
/////////////////////////////////////////////////////////////////////////////////

module pdec_reg_dyn_bd (
    //System
    input               rst_n            ,
    input               clk              ,

    //w/r interface
    input               wen              ,
    input               ren              ,
    input      [32-1:0] waddr            ,
    input      [32-1:0] raddr            ,
    input      [32-1:0] wdata            ,
    output reg [32-1:0] rdata            ,

    //common_para
    output reg [ 2-1:0] dcrc_num         ,
    output reg [ 2-1:0] list_num         ,
    output reg          leaf_mode        ,
    output reg [ 9-1:0] param_k          ,
    output reg [ 9-1:0] param_a          ,
    output reg [ 3-1:0] param_n          ,

    //jump_type0
    output reg [32-1:0] jump_type0       ,

    //jump_type1
    output reg [32-1:0] jump_type1       ,

    //jump_type2
    output reg [32-1:0] jump_type2       ,

    //jump_type3
    output reg [32-1:0] jump_type3       ,

    //jump_type4
    output reg [32-1:0] jump_type4       ,

    //jump_type5
    output reg [32-1:0] jump_type5       ,

    //jump_type6
    output reg [32-1:0] jump_type6       ,

    //jump_type7
    output reg [32-1:0] jump_type7       ,

    //jump_type8
    output reg [32-1:0] jump_type8       ,

    //jump_type9
    output reg [32-1:0] jump_type9       ,

    //jump_type10
    output reg [32-1:0] jump_type10      ,

    //jump_type11
    output reg [32-1:0] jump_type11      ,

    //jump_type12
    output reg [32-1:0] jump_type12      ,

    //jump_type13
    output reg [32-1:0] jump_type13      ,

    //jump_type14
    output reg [32-1:0] jump_type14      ,

    //jump_type15
    output reg [32-1:0] jump_type15      ,

    //jump_type16
    output reg [32-1:0] jump_type16      ,

    //jump_type17
    output reg [32-1:0] jump_type17      ,

    //jump_type18
    output reg [32-1:0] jump_type18      ,

    //jump_type19
    output reg [32-1:0] jump_type19      ,

    //jump_type20
    output reg [32-1:0] jump_type20      ,

    //jump_type21
    output reg [32-1:0] jump_type21      ,

    //jump_type22
    output reg [32-1:0] jump_type22      ,

    //jump_type23
    output reg [32-1:0] jump_type23      ,

    //jump_type24
    output reg [32-1:0] jump_type24      ,

    //jump_type25
    output reg [32-1:0] jump_type25      ,

    //jump_type26
    output reg [32-1:0] jump_type26      ,

    //jump_type27
    output reg [32-1:0] jump_type27      ,

    //jump_type28
    output reg [32-1:0] jump_type28      ,

    //jump_type29
    output reg [32-1:0] jump_type29      ,

    //jump_type30
    output reg [32-1:0] jump_type30      ,

    //jump_type31
    output reg [32-1:0] jump_type31      ,

    //jump_type32
    output reg [32-1:0] jump_type32      ,

    //jump_type33
    output reg [32-1:0] jump_type33      ,

    //jump_type34
    output reg [32-1:0] jump_type34      ,

    //jump_type35
    output reg [32-1:0] jump_type35      ,

    //jump_type36
    output reg [32-1:0] jump_type36      ,

    //jump_type37
    output reg [32-1:0] jump_type37      ,

    //jump_type38
    output reg [32-1:0] jump_type38      ,

    //jump_type39
    output reg [32-1:0] jump_type39      ,

    //jump_type40
    output reg [32-1:0] jump_type40      ,

    //jump_type41
    output reg [32-1:0] jump_type41      ,

    //jump_type42
    output reg [32-1:0] jump_type42      ,

    //jump_type43
    output reg [32-1:0] jump_type43      ,

    //jump_type44
    output reg [32-1:0] jump_type44      ,

    //jump_type45
    output reg [32-1:0] jump_type45      ,

    //jump_type46
    output reg [32-1:0] jump_type46      ,

    //jump_type47
    output reg [32-1:0] jump_type47      ,

    //jump_type48
    output reg [32-1:0] jump_type48      ,

    //jump_type49
    output reg [32-1:0] jump_type49      ,

    //jump_type50
    output reg [32-1:0] jump_type50      ,

    //jump_type51
    output reg [32-1:0] jump_type51      ,

    //jump_type52
    output reg [32-1:0] jump_type52      ,

    //jump_type53
    output reg [32-1:0] jump_type53      ,

    //jump_type54
    output reg [32-1:0] jump_type54      ,

    //jump_type55
    output reg [32-1:0] jump_type55      ,

    //jump_type56
    output reg [32-1:0] jump_type56      ,

    //jump_type57
    output reg [32-1:0] jump_type57      ,

    //jump_type58
    output reg [32-1:0] jump_type58      ,

    //jump_type59
    output reg [32-1:0] jump_type59      ,

    //jump_type60
    output reg [32-1:0] jump_type60      ,

    //jump_type61
    output reg [32-1:0] jump_type61      ,

    //jump_type62
    output reg [32-1:0] jump_type62      ,

    //jump_type63
    output reg [32-1:0] jump_type63      ,

    //jump_type64
    output reg [32-1:0] jump_type64      ,

    //jump_type65
    output reg [32-1:0] jump_type65      ,

    //jump_type66
    output reg [32-1:0] jump_type66      ,

    //jump_type67
    output reg [32-1:0] jump_type67      ,

    //jump_type68
    output reg [32-1:0] jump_type68      ,

    //jump_type69
    output reg [32-1:0] jump_type69      ,

    //jump_type70
    output reg [32-1:0] jump_type70      ,

    //jump_type71
    output reg [32-1:0] jump_type71      ,

    //jump_type72
    output reg [32-1:0] jump_type72      ,

    //jump_type73
    output reg [32-1:0] jump_type73      ,

    //jump_type74
    output reg [32-1:0] jump_type74      ,

    //jump_type75
    output reg [32-1:0] jump_type75      ,

    //jump_type76
    output reg [32-1:0] jump_type76      ,

    //jump_type77
    output reg [32-1:0] jump_type77      ,

    //jump_type78
    output reg [32-1:0] jump_type78      ,

    //jump_type79
    output reg [32-1:0] jump_type79      ,

    //jump_type80
    output reg [32-1:0] jump_type80      ,

    //jump_type81
    output reg [32-1:0] jump_type81      ,

    //jump_type82
    output reg [32-1:0] jump_type82      ,

    //jump_type83
    output reg [32-1:0] jump_type83      ,

    //jump_type84
    output reg [32-1:0] jump_type84      ,

    //jump_type85
    output reg [32-1:0] jump_type85      ,

    //jump_type86
    output reg [32-1:0] jump_type86      ,

    //jump_type87
    output reg [32-1:0] jump_type87      ,

    //jump_type88
    output reg [32-1:0] jump_type88      ,

    //jump_type89
    output reg [32-1:0] jump_type89      ,

    //jump_type90
    output reg [32-1:0] jump_type90      ,

    //jump_type91
    output reg [32-1:0] jump_type91      ,

    //jump_type92
    output reg [32-1:0] jump_type92      ,

    //jump_type93
    output reg [32-1:0] jump_type93      ,

    //jump_type94
    output reg [32-1:0] jump_type94      ,

    //jump_type95
    output reg [32-1:0] jump_type95      ,

    //jump_type96
    output reg [32-1:0] jump_type96      ,

    //jump_type97
    output reg [32-1:0] jump_type97      ,

    //jump_type98
    output reg [32-1:0] jump_type98      ,

    //jump_type99
    output reg [32-1:0] jump_type99      ,

    //jump_type100
    output reg [32-1:0] jump_type100     ,

    //jump_type101
    output reg [32-1:0] jump_type101     ,

    //jump_type102
    output reg [32-1:0] jump_type102     ,

    //jump_type103
    output reg [32-1:0] jump_type103     ,

    //jump_type104
    output reg [32-1:0] jump_type104     ,

    //jump_type105
    output reg [32-1:0] jump_type105     ,

    //jump_type106
    output reg [32-1:0] jump_type106     ,

    //jump_type107
    output reg [32-1:0] jump_type107     ,

    //jump_type108
    output reg [32-1:0] jump_type108     ,

    //jump_type109
    output reg [32-1:0] jump_type109     ,

    //jump_type110
    output reg [32-1:0] jump_type110     ,

    //jump_type111
    output reg [32-1:0] jump_type111     ,

    //jump_type112
    output reg [32-1:0] jump_type112     ,

    //jump_type113
    output reg [32-1:0] jump_type113     ,

    //jump_type114
    output reg [32-1:0] jump_type114     ,

    //jump_type115
    output reg [32-1:0] jump_type115     ,

    //jump_type116
    output reg [32-1:0] jump_type116     ,

    //jump_type117
    output reg [32-1:0] jump_type117     ,

    //jump_type118
    output reg [32-1:0] jump_type118     ,

    //jump_type119
    output reg [32-1:0] jump_type119     ,

    //jump_type120
    output reg [32-1:0] jump_type120     ,

    //jump_type121
    output reg [32-1:0] jump_type121     ,

    //jump_type122
    output reg [32-1:0] jump_type122     ,

    //jump_type123
    output reg [32-1:0] jump_type123     ,

    //jump_type124
    output reg [32-1:0] jump_type124     ,

    //jump_type125
    output reg [32-1:0] jump_type125     ,

    //jump_type126
    output reg [32-1:0] jump_type126     ,

    //jump_type127
    output reg [32-1:0] jump_type127     ,

    //jump_type128
    output reg [32-1:0] jump_type128     ,

    //jump_type129
    output reg [32-1:0] jump_type129     ,

    //jump_type130
    output reg [32-1:0] jump_type130     ,

    //jump_type131
    output reg [32-1:0] jump_type131     ,

    //jump_type132
    output reg [32-1:0] jump_type132     ,

    //jump_type133
    output reg [32-1:0] jump_type133     ,

    //jump_type134
    output reg [32-1:0] jump_type134     ,

    //jump_type135
    output reg [32-1:0] jump_type135     ,

    //jump_type136
    output reg [32-1:0] jump_type136     ,

    //jump_type137
    output reg [32-1:0] jump_type137     ,

    //jump_type138
    output reg [32-1:0] jump_type138     ,

    //jump_type139
    output reg [32-1:0] jump_type139     ,

    //jump_type140
    output reg [32-1:0] jump_type140     ,

    //jump_type141
    output reg [32-1:0] jump_type141     ,

    //jump_type142
    output reg [32-1:0] jump_type142     ,

    //jump_type143
    output reg [32-1:0] jump_type143     ,

    //jump_type144
    output reg [32-1:0] jump_type144     ,

    //jump_type145
    output reg [32-1:0] jump_type145     ,

    //jump_type146
    output reg [32-1:0] jump_type146     ,

    //jump_type147
    output reg [32-1:0] jump_type147     ,

    //jump_type148
    output reg [32-1:0] jump_type148     ,

    //jump_type149
    output reg [32-1:0] jump_type149     ,

    //jump_type150
    output reg [32-1:0] jump_type150     ,

    //jump_type151
    output reg [32-1:0] jump_type151     ,

    //jump_type152
    output reg [32-1:0] jump_type152     ,

    //jump_type153
    output reg [32-1:0] jump_type153     ,

    //jump_type154
    output reg [32-1:0] jump_type154     ,

    //jump_type155
    output reg [32-1:0] jump_type155     ,

    //jump_type156
    output reg [32-1:0] jump_type156     ,

    //jump_type157
    output reg [32-1:0] jump_type157     ,

    //jump_type158
    output reg [32-1:0] jump_type158     ,

    //jump_type159
    output reg [32-1:0] jump_type159     ,

    //jump_type160
    output reg [32-1:0] jump_type160     ,

    //jump_type161
    output reg [32-1:0] jump_type161     ,

    //jump_type162
    output reg [32-1:0] jump_type162     ,

    //jump_type163
    output reg [32-1:0] jump_type163     ,

    //jump_type164
    output reg [32-1:0] jump_type164     ,

    //jump_type165
    output reg [32-1:0] jump_type165     ,

    //jump_type166
    output reg [32-1:0] jump_type166     ,

    //jump_type167
    output reg [32-1:0] jump_type167     ,

    //jump_type168
    output reg [32-1:0] jump_type168     ,

    //jump_type169
    output reg [32-1:0] jump_type169     ,

    //jump_type170
    output reg [32-1:0] jump_type170     ,

    //jump_type171
    output reg [32-1:0] jump_type171     ,

    //jump_type172
    output reg [32-1:0] jump_type172     ,

    //jump_type173
    output reg [32-1:0] jump_type173     ,

    //jump_type174
    output reg [32-1:0] jump_type174     ,

    //jump_type175
    output reg [32-1:0] jump_type175     ,

    //jump_type176
    output reg [32-1:0] jump_type176     ,

    //jump_type177
    output reg [32-1:0] jump_type177     ,

    //jump_type178
    output reg [32-1:0] jump_type178     ,

    //jump_type179
    output reg [32-1:0] jump_type179     ,

    //jump_type180
    output reg [32-1:0] jump_type180     ,

    //jump_type181
    output reg [32-1:0] jump_type181     ,

    //jump_type182
    output reg [32-1:0] jump_type182     ,

    //jump_type183
    output reg [32-1:0] jump_type183     ,

    //jump_type184
    output reg [32-1:0] jump_type184     ,

    //jump_type185
    output reg [32-1:0] jump_type185     ,

    //jump_type186
    output reg [32-1:0] jump_type186     ,

    //jump_type187
    output reg [32-1:0] jump_type187     ,

    //jump_type188
    output reg [32-1:0] jump_type188     ,

    //jump_type189
    output reg [32-1:0] jump_type189     ,

    //jump_type190
    output reg [32-1:0] jump_type190     ,

    //jump_type191
    output reg [32-1:0] jump_type191     ,

    //jump_type192
    output reg [32-1:0] jump_type192     ,

    //jump_type193
    output reg [32-1:0] jump_type193     ,

    //jump_type194
    output reg [32-1:0] jump_type194     ,

    //jump_type195
    output reg [32-1:0] jump_type195     ,

    //jump_type196
    output reg [32-1:0] jump_type196     ,

    //jump_type197
    output reg [32-1:0] jump_type197     ,

    //jump_type198
    output reg [32-1:0] jump_type198     ,

    //jump_type199
    output reg [32-1:0] jump_type199     ,

    //jump_type200
    output reg [32-1:0] jump_type200     ,

    //jump_type201
    output reg [32-1:0] jump_type201     ,

    //jump_type202
    output reg [32-1:0] jump_type202     ,

    //jump_type203
    output reg [32-1:0] jump_type203     ,

    //jump_type204
    output reg [32-1:0] jump_type204     ,

    //jump_type205
    output reg [32-1:0] jump_type205     ,

    //jump_type206
    output reg [32-1:0] jump_type206     ,

    //jump_type207
    output reg [32-1:0] jump_type207     ,

    //jump_type208
    output reg [32-1:0] jump_type208     ,

    //jump_type209
    output reg [32-1:0] jump_type209     ,

    //jump_type210
    output reg [32-1:0] jump_type210     ,

    //jump_type211
    output reg [32-1:0] jump_type211     ,

    //jump_type212
    output reg [32-1:0] jump_type212     ,

    //jump_type213
    output reg [32-1:0] jump_type213     ,

    //jump_type214
    output reg [32-1:0] jump_type214     ,

    //jump_type215
    output reg [32-1:0] jump_type215     ,

    //jump_type216
    output reg [32-1:0] jump_type216     ,

    //jump_type217
    output reg [32-1:0] jump_type217     ,

    //jump_type218
    output reg [32-1:0] jump_type218     ,

    //jump_type219
    output reg [32-1:0] jump_type219     ,

    //jump_type220
    output reg [32-1:0] jump_type220     ,

    //jump_type221
    output reg [32-1:0] jump_type221     ,

    //jump_type222
    output reg [32-1:0] jump_type222     ,

    //jump_type223
    output reg [32-1:0] jump_type223     ,

    //jump_type224
    output reg [32-1:0] jump_type224     ,

    //jump_type225
    output reg [32-1:0] jump_type225     ,

    //jump_type226
    output reg [32-1:0] jump_type226     ,

    //jump_type227
    output reg [32-1:0] jump_type227     ,

    //jump_type228
    output reg [32-1:0] jump_type228     ,

    //jump_type229
    output reg [32-1:0] jump_type229     ,

    //jump_type230
    output reg [32-1:0] jump_type230     ,

    //jump_type231
    output reg [32-1:0] jump_type231     ,

    //jump_type232
    output reg [32-1:0] jump_type232     ,

    //jump_type233
    output reg [32-1:0] jump_type233     ,

    //jump_type234
    output reg [32-1:0] jump_type234     ,

    //jump_type235
    output reg [32-1:0] jump_type235     ,

    //jump_type236
    output reg [32-1:0] jump_type236     ,

    //jump_type237
    output reg [32-1:0] jump_type237     ,

    //jump_type238
    output reg [32-1:0] jump_type238     ,

    //jump_type239
    output reg [32-1:0] jump_type239     ,

    //jump_type240
    output reg [32-1:0] jump_type240     ,

    //jump_type241
    output reg [32-1:0] jump_type241     ,

    //jump_type242
    output reg [32-1:0] jump_type242     ,

    //jump_type243
    output reg [32-1:0] jump_type243     ,

    //jump_type244
    output reg [32-1:0] jump_type244     ,

    //jump_type245
    output reg [32-1:0] jump_type245     ,

    //jump_type246
    output reg [32-1:0] jump_type246     ,

    //jump_type247
    output reg [32-1:0] jump_type247     ,

    //jump_type248
    output reg [32-1:0] jump_type248     ,

    //jump_type249
    output reg [32-1:0] jump_type249     ,

    //jump_type250
    output reg [32-1:0] jump_type250     ,

    //jump_type251
    output reg [32-1:0] jump_type251     ,

    //jump_type252
    output reg [32-1:0] jump_type252     ,

    //jump_type253
    output reg [32-1:0] jump_type253     ,

    //jump_type254
    output reg [32-1:0] jump_type254     ,

    //jump_type255
    output reg [32-1:0] jump_type255     ,

    //jump_type256
    output reg [32-1:0] jump_type256     ,

    //jump_type257
    output reg [32-1:0] jump_type257     ,

    //jump_type258
    output reg [32-1:0] jump_type258     ,

    //jump_type259
    output reg [32-1:0] jump_type259     ,

    //jump_type260
    output reg [32-1:0] jump_type260     ,

    //jump_type261
    output reg [32-1:0] jump_type261     ,

    //jump_type262
    output reg [32-1:0] jump_type262     ,

    //jump_type263
    output reg [32-1:0] jump_type263     ,

    //jump_type264
    output reg [32-1:0] jump_type264     ,

    //jump_type265
    output reg [32-1:0] jump_type265     ,

    //jump_type266
    output reg [32-1:0] jump_type266     ,

    //jump_type267
    output reg [32-1:0] jump_type267     ,

    //jump_type268
    output reg [32-1:0] jump_type268     ,

    //jump_type269
    output reg [32-1:0] jump_type269     ,

    //jump_type270
    output reg [32-1:0] jump_type270     ,

    //jump_type271
    output reg [32-1:0] jump_type271     ,

    //jump_type272
    output reg [32-1:0] jump_type272     ,

    //jump_type273
    output reg [32-1:0] jump_type273     ,

    //jump_type274
    output reg [32-1:0] jump_type274     ,

    //jump_type275
    output reg [32-1:0] jump_type275     ,

    //jump_type276
    output reg [32-1:0] jump_type276     ,

    //jump_type277
    output reg [32-1:0] jump_type277     ,

    //jump_type278
    output reg [32-1:0] jump_type278     ,

    //jump_type279
    output reg [32-1:0] jump_type279     ,

    //jump_type280
    output reg [32-1:0] jump_type280     ,

    //jump_type281
    output reg [32-1:0] jump_type281     ,

    //jump_type282
    output reg [32-1:0] jump_type282     ,

    //jump_type283
    output reg [32-1:0] jump_type283     ,

    //jump_type284
    output reg [32-1:0] jump_type284     ,

    //jump_type285
    output reg [32-1:0] jump_type285     ,

    //jump_type286
    output reg [32-1:0] jump_type286     ,

    //jump_type287
    output reg [32-1:0] jump_type287     ,

    //jump_type288
    output reg [32-1:0] jump_type288     ,

    //jump_type289
    output reg [32-1:0] jump_type289     ,

    //jump_type290
    output reg [32-1:0] jump_type290     ,

    //jump_type291
    output reg [32-1:0] jump_type291     ,

    //jump_type292
    output reg [32-1:0] jump_type292     ,

    //jump_type293
    output reg [32-1:0] jump_type293     ,

    //jump_type294
    output reg [32-1:0] jump_type294     ,

    //jump_type295
    output reg [32-1:0] jump_type295     ,

    //jump_type296
    output reg [32-1:0] jump_type296     ,

    //jump_type297
    output reg [32-1:0] jump_type297     ,

    //jump_type298
    output reg [32-1:0] jump_type298     ,

    //jump_type299
    output reg [32-1:0] jump_type299     ,

    //jump_type300
    output reg [32-1:0] jump_type300     ,

    //jump_type301
    output reg [32-1:0] jump_type301     ,

    //jump_type302
    output reg [32-1:0] jump_type302     ,

    //jump_type303
    output reg [32-1:0] jump_type303     ,

    //jump_type304
    output reg [32-1:0] jump_type304     ,

    //jump_type305
    output reg [32-1:0] jump_type305     ,

    //jump_type306
    output reg [32-1:0] jump_type306     ,

    //jump_type307
    output reg [32-1:0] jump_type307     ,

    //jump_type308
    output reg [32-1:0] jump_type308     ,

    //jump_type309
    output reg [32-1:0] jump_type309     ,

    //jump_type310
    output reg [32-1:0] jump_type310     ,

    //jump_type311
    output reg [32-1:0] jump_type311     ,

    //jump_type312
    output reg [32-1:0] jump_type312     ,

    //jump_type313
    output reg [32-1:0] jump_type313     ,

    //jump_type314
    output reg [32-1:0] jump_type314     ,

    //jump_type315
    output reg [32-1:0] jump_type315     ,

    //jump_type316
    output reg [32-1:0] jump_type316     ,

    //jump_type317
    output reg [32-1:0] jump_type317     ,

    //jump_type318
    output reg [32-1:0] jump_type318     ,

    //jump_type319
    output reg [32-1:0] jump_type319     ,

    //jump_type320
    output reg [32-1:0] jump_type320     ,

    //jump_type321
    output reg [32-1:0] jump_type321     ,

    //jump_type322
    output reg [32-1:0] jump_type322     ,

    //jump_type323
    output reg [32-1:0] jump_type323     ,

    //jump_type324
    output reg [32-1:0] jump_type324     ,

    //jump_type325
    output reg [32-1:0] jump_type325     ,

    //jump_type326
    output reg [32-1:0] jump_type326     ,

    //jump_type327
    output reg [32-1:0] jump_type327     ,

    //jump_type328
    output reg [32-1:0] jump_type328     ,

    //jump_type329
    output reg [32-1:0] jump_type329     ,

    //jump_type330
    output reg [32-1:0] jump_type330     ,

    //jump_type331
    output reg [32-1:0] jump_type331     ,

    //jump_type332
    output reg [32-1:0] jump_type332     ,

    //jump_type333
    output reg [32-1:0] jump_type333     ,

    //jump_type334
    output reg [32-1:0] jump_type334     ,

    //jump_type335
    output reg [32-1:0] jump_type335     ,

    //jump_type336
    output reg [32-1:0] jump_type336     ,

    //jump_type337
    output reg [32-1:0] jump_type337     ,

    //jump_type338
    output reg [32-1:0] jump_type338     ,

    //jump_type339
    output reg [32-1:0] jump_type339     ,

    //jump_type340
    output reg [32-1:0] jump_type340     ,

    //jump_type341
    output reg [32-1:0] jump_type341     ,

    //jump_type342
    output reg [32-1:0] jump_type342     ,

    //jump_type343
    output reg [32-1:0] jump_type343     ,

    //jump_type344
    output reg [32-1:0] jump_type344     ,

    //jump_type345
    output reg [32-1:0] jump_type345     ,

    //jump_type346
    output reg [32-1:0] jump_type346     ,

    //jump_type347
    output reg [32-1:0] jump_type347     ,

    //jump_type348
    output reg [32-1:0] jump_type348     ,

    //jump_type349
    output reg [32-1:0] jump_type349     ,

    //jump_type350
    output reg [32-1:0] jump_type350     ,

    //jump_type351
    output reg [32-1:0] jump_type351     ,

    //jump_type352
    output reg [32-1:0] jump_type352     ,

    //jump_type353
    output reg [32-1:0] jump_type353     ,

    //jump_type354
    output reg [32-1:0] jump_type354     ,

    //jump_type355
    output reg [32-1:0] jump_type355     ,

    //jump_type356
    output reg [32-1:0] jump_type356     ,

    //jump_type357
    output reg [32-1:0] jump_type357     ,

    //jump_type358
    output reg [32-1:0] jump_type358     ,

    //jump_type359
    output reg [32-1:0] jump_type359     ,

    //jump_type360
    output reg [32-1:0] jump_type360     ,

    //jump_type361
    output reg [32-1:0] jump_type361     ,

    //jump_type362
    output reg [32-1:0] jump_type362     ,

    //jump_type363
    output reg [32-1:0] jump_type363     ,

    //jump_type364
    output reg [32-1:0] jump_type364     ,

    //jump_type365
    output reg [32-1:0] jump_type365     ,

    //jump_type366
    output reg [32-1:0] jump_type366     ,

    //jump_type367
    output reg [32-1:0] jump_type367     ,

    //jump_type368
    output reg [32-1:0] jump_type368     ,

    //jump_type369
    output reg [32-1:0] jump_type369     ,

    //jump_type370
    output reg [32-1:0] jump_type370     ,

    //jump_type371
    output reg [32-1:0] jump_type371     ,

    //jump_type372
    output reg [32-1:0] jump_type372     ,

    //jump_type373
    output reg [32-1:0] jump_type373     ,

    //jump_type374
    output reg [32-1:0] jump_type374     ,

    //jump_type375
    output reg [32-1:0] jump_type375     ,

    //jump_type376
    output reg [32-1:0] jump_type376     ,

    //jump_type377
    output reg [32-1:0] jump_type377     ,

    //jump_type378
    output reg [32-1:0] jump_type378     ,

    //jump_type379
    output reg [32-1:0] jump_type379     ,

    //jump_type380
    output reg [32-1:0] jump_type380     ,

    //jump_type381
    output reg [32-1:0] jump_type381     ,

    //jump_type382
    output reg [32-1:0] jump_type382     ,

    //jump_type383
    output reg [32-1:0] jump_type383     ,

    //jump_type384
    output reg [32-1:0] jump_type384     ,

    //jump_type385
    output reg [32-1:0] jump_type385     ,

    //jump_type386
    output reg [32-1:0] jump_type386     ,

    //jump_type387
    output reg [32-1:0] jump_type387     ,

    //jump_type388
    output reg [32-1:0] jump_type388     ,

    //jump_type389
    output reg [32-1:0] jump_type389     ,

    //jump_type390
    output reg [32-1:0] jump_type390     ,

    //jump_type391
    output reg [32-1:0] jump_type391     ,

    //jump_type392
    output reg [32-1:0] jump_type392     ,

    //jump_type393
    output reg [32-1:0] jump_type393     ,

    //jump_type394
    output reg [32-1:0] jump_type394     ,

    //jump_type395
    output reg [32-1:0] jump_type395     ,

    //jump_type396
    output reg [32-1:0] jump_type396     ,

    //jump_type397
    output reg [32-1:0] jump_type397     ,

    //jump_type398
    output reg [32-1:0] jump_type398     ,

    //jump_type399
    output reg [32-1:0] jump_type399     ,

    //jump_type400
    output reg [32-1:0] jump_type400     ,

    //jump_type401
    output reg [32-1:0] jump_type401     ,

    //jump_type402
    output reg [32-1:0] jump_type402     ,

    //jump_type403
    output reg [32-1:0] jump_type403     ,

    //jump_type404
    output reg [32-1:0] jump_type404     ,

    //jump_type405
    output reg [32-1:0] jump_type405     ,

    //jump_type406
    output reg [32-1:0] jump_type406     ,

    //jump_type407
    output reg [32-1:0] jump_type407     ,

    //jump_type408
    output reg [32-1:0] jump_type408     ,

    //jump_type409
    output reg [32-1:0] jump_type409     ,

    //jump_type410
    output reg [32-1:0] jump_type410     ,

    //jump_type411
    output reg [32-1:0] jump_type411     ,

    //jump_type412
    output reg [32-1:0] jump_type412     ,

    //jump_type413
    output reg [32-1:0] jump_type413     ,

    //jump_type414
    output reg [32-1:0] jump_type414     ,

    //jump_type415
    output reg [32-1:0] jump_type415     ,

    //jump_type416
    output reg [32-1:0] jump_type416     ,

    //jump_type417
    output reg [32-1:0] jump_type417     ,

    //jump_type418
    output reg [32-1:0] jump_type418     ,

    //jump_type419
    output reg [32-1:0] jump_type419     ,

    //jump_type420
    output reg [32-1:0] jump_type420     ,

    //jump_type421
    output reg [32-1:0] jump_type421     ,

    //jump_type422
    output reg [32-1:0] jump_type422     ,

    //jump_type423
    output reg [32-1:0] jump_type423     ,

    //jump_type424
    output reg [32-1:0] jump_type424     ,

    //jump_type425
    output reg [32-1:0] jump_type425     ,

    //jump_type426
    output reg [32-1:0] jump_type426     ,

    //jump_type427
    output reg [32-1:0] jump_type427     ,

    //jump_type428
    output reg [32-1:0] jump_type428     ,

    //jump_type429
    output reg [32-1:0] jump_type429     ,

    //jump_type430
    output reg [32-1:0] jump_type430     ,

    //jump_type431
    output reg [32-1:0] jump_type431     ,

    //jump_type432
    output reg [32-1:0] jump_type432     ,

    //jump_type433
    output reg [32-1:0] jump_type433     ,

    //jump_type434
    output reg [32-1:0] jump_type434     ,

    //jump_type435
    output reg [32-1:0] jump_type435     ,

    //jump_type436
    output reg [32-1:0] jump_type436     ,

    //jump_type437
    output reg [32-1:0] jump_type437     ,

    //jump_type438
    output reg [32-1:0] jump_type438     ,

    //jump_type439
    output reg [32-1:0] jump_type439     ,

    //jump_type440
    output reg [32-1:0] jump_type440     ,

    //jump_type441
    output reg [32-1:0] jump_type441     ,

    //jump_type442
    output reg [32-1:0] jump_type442     ,

    //jump_type443
    output reg [32-1:0] jump_type443     ,

    //jump_type444
    output reg [32-1:0] jump_type444     ,

    //jump_type445
    output reg [32-1:0] jump_type445     ,

    //jump_type446
    output reg [32-1:0] jump_type446     ,

    //jump_type447
    output reg [32-1:0] jump_type447     ,

    //jump_type448
    output reg [32-1:0] jump_type448     ,

    //jump_type449
    output reg [32-1:0] jump_type449     ,

    //jump_type450
    output reg [32-1:0] jump_type450     ,

    //jump_type451
    output reg [32-1:0] jump_type451     ,

    //jump_type452
    output reg [32-1:0] jump_type452     ,

    //jump_type453
    output reg [32-1:0] jump_type453     ,

    //jump_type454
    output reg [32-1:0] jump_type454     ,

    //jump_type455
    output reg [32-1:0] jump_type455     ,

    //jump_type456
    output reg [32-1:0] jump_type456     ,

    //jump_type457
    output reg [32-1:0] jump_type457     ,

    //jump_type458
    output reg [32-1:0] jump_type458     ,

    //jump_type459
    output reg [32-1:0] jump_type459     ,

    //jump_type460
    output reg [32-1:0] jump_type460     ,

    //jump_type461
    output reg [32-1:0] jump_type461     ,

    //jump_type462
    output reg [32-1:0] jump_type462     ,

    //jump_type463
    output reg [32-1:0] jump_type463     ,

    //jump_type464
    output reg [32-1:0] jump_type464     ,

    //jump_type465
    output reg [32-1:0] jump_type465     ,

    //jump_type466
    output reg [32-1:0] jump_type466     ,

    //jump_type467
    output reg [32-1:0] jump_type467     ,

    //jump_type468
    output reg [32-1:0] jump_type468     ,

    //jump_type469
    output reg [32-1:0] jump_type469     ,

    //jump_type470
    output reg [32-1:0] jump_type470     ,

    //jump_type471
    output reg [32-1:0] jump_type471     ,

    //jump_type472
    output reg [32-1:0] jump_type472     ,

    //jump_type473
    output reg [32-1:0] jump_type473     ,

    //jump_type474
    output reg [32-1:0] jump_type474     ,

    //jump_type475
    output reg [32-1:0] jump_type475     ,

    //jump_type476
    output reg [32-1:0] jump_type476     ,

    //jump_type477
    output reg [32-1:0] jump_type477     ,

    //jump_type478
    output reg [32-1:0] jump_type478     ,

    //jump_type479
    output reg [32-1:0] jump_type479     ,

    //jump_type480
    output reg [32-1:0] jump_type480     ,

    //jump_type481
    output reg [32-1:0] jump_type481     ,

    //jump_type482
    output reg [32-1:0] jump_type482     ,

    //jump_type483
    output reg [32-1:0] jump_type483     ,

    //jump_type484
    output reg [32-1:0] jump_type484     ,

    //jump_type485
    output reg [32-1:0] jump_type485     ,

    //jump_type486
    output reg [32-1:0] jump_type486     ,

    //jump_type487
    output reg [32-1:0] jump_type487     ,

    //jump_type488
    output reg [32-1:0] jump_type488     ,

    //jump_type489
    output reg [32-1:0] jump_type489     ,

    //jump_type490
    output reg [32-1:0] jump_type490     ,

    //jump_type491
    output reg [32-1:0] jump_type491     ,

    //jump_type492
    output reg [32-1:0] jump_type492     ,

    //jump_type493
    output reg [32-1:0] jump_type493     ,

    //jump_type494
    output reg [32-1:0] jump_type494     ,

    //jump_type495
    output reg [32-1:0] jump_type495     ,

    //jump_type496
    output reg [32-1:0] jump_type496     ,

    //jump_type497
    output reg [32-1:0] jump_type497     ,

    //jump_type498
    output reg [32-1:0] jump_type498     ,

    //jump_type499
    output reg [32-1:0] jump_type499     ,

    //jump_type500
    output reg [32-1:0] jump_type500     ,

    //jump_type501
    output reg [32-1:0] jump_type501     ,

    //jump_type502
    output reg [32-1:0] jump_type502     ,

    //jump_type503
    output reg [32-1:0] jump_type503     ,

    //jump_type504
    output reg [32-1:0] jump_type504     ,

    //jump_type505
    output reg [32-1:0] jump_type505     ,

    //jump_type506
    output reg [32-1:0] jump_type506     ,

    //jump_type507
    output reg [32-1:0] jump_type507     ,

    //jump_type508
    output reg [32-1:0] jump_type508     ,

    //jump_type509
    output reg [32-1:0] jump_type509     ,

    //jump_type510
    output reg [32-1:0] jump_type510     ,

    //jump_type511
    output reg [28-1:0] jump_type511     
);

//----------------------------local parameter---------------------------------------------
localparam COMMON_PARA_REG          = 32'h0  ;
localparam JUMP_TYPE0_REG           = 32'h4  ;
localparam JUMP_TYPE1_REG           = 32'h8  ;
localparam JUMP_TYPE2_REG           = 32'hc  ;
localparam JUMP_TYPE3_REG           = 32'h10 ;
localparam JUMP_TYPE4_REG           = 32'h14 ;
localparam JUMP_TYPE5_REG           = 32'h18 ;
localparam JUMP_TYPE6_REG           = 32'h1c ;
localparam JUMP_TYPE7_REG           = 32'h20 ;
localparam JUMP_TYPE8_REG           = 32'h24 ;
localparam JUMP_TYPE9_REG           = 32'h28 ;
localparam JUMP_TYPE10_REG          = 32'h2c ;
localparam JUMP_TYPE11_REG          = 32'h30 ;
localparam JUMP_TYPE12_REG          = 32'h34 ;
localparam JUMP_TYPE13_REG          = 32'h38 ;
localparam JUMP_TYPE14_REG          = 32'h3c ;
localparam JUMP_TYPE15_REG          = 32'h40 ;
localparam JUMP_TYPE16_REG          = 32'h44 ;
localparam JUMP_TYPE17_REG          = 32'h48 ;
localparam JUMP_TYPE18_REG          = 32'h4c ;
localparam JUMP_TYPE19_REG          = 32'h50 ;
localparam JUMP_TYPE20_REG          = 32'h54 ;
localparam JUMP_TYPE21_REG          = 32'h58 ;
localparam JUMP_TYPE22_REG          = 32'h5c ;
localparam JUMP_TYPE23_REG          = 32'h60 ;
localparam JUMP_TYPE24_REG          = 32'h64 ;
localparam JUMP_TYPE25_REG          = 32'h68 ;
localparam JUMP_TYPE26_REG          = 32'h6c ;
localparam JUMP_TYPE27_REG          = 32'h70 ;
localparam JUMP_TYPE28_REG          = 32'h74 ;
localparam JUMP_TYPE29_REG          = 32'h78 ;
localparam JUMP_TYPE30_REG          = 32'h7c ;
localparam JUMP_TYPE31_REG          = 32'h80 ;
localparam JUMP_TYPE32_REG          = 32'h84 ;
localparam JUMP_TYPE33_REG          = 32'h88 ;
localparam JUMP_TYPE34_REG          = 32'h8c ;
localparam JUMP_TYPE35_REG          = 32'h90 ;
localparam JUMP_TYPE36_REG          = 32'h94 ;
localparam JUMP_TYPE37_REG          = 32'h98 ;
localparam JUMP_TYPE38_REG          = 32'h9c ;
localparam JUMP_TYPE39_REG          = 32'ha0 ;
localparam JUMP_TYPE40_REG          = 32'ha4 ;
localparam JUMP_TYPE41_REG          = 32'ha8 ;
localparam JUMP_TYPE42_REG          = 32'hac ;
localparam JUMP_TYPE43_REG          = 32'hb0 ;
localparam JUMP_TYPE44_REG          = 32'hb4 ;
localparam JUMP_TYPE45_REG          = 32'hb8 ;
localparam JUMP_TYPE46_REG          = 32'hbc ;
localparam JUMP_TYPE47_REG          = 32'hc0 ;
localparam JUMP_TYPE48_REG          = 32'hc4 ;
localparam JUMP_TYPE49_REG          = 32'hc8 ;
localparam JUMP_TYPE50_REG          = 32'hcc ;
localparam JUMP_TYPE51_REG          = 32'hd0 ;
localparam JUMP_TYPE52_REG          = 32'hd4 ;
localparam JUMP_TYPE53_REG          = 32'hd8 ;
localparam JUMP_TYPE54_REG          = 32'hdc ;
localparam JUMP_TYPE55_REG          = 32'he0 ;
localparam JUMP_TYPE56_REG          = 32'he4 ;
localparam JUMP_TYPE57_REG          = 32'he8 ;
localparam JUMP_TYPE58_REG          = 32'hec ;
localparam JUMP_TYPE59_REG          = 32'hf0 ;
localparam JUMP_TYPE60_REG          = 32'hf4 ;
localparam JUMP_TYPE61_REG          = 32'hf8 ;
localparam JUMP_TYPE62_REG          = 32'hfc ;
localparam JUMP_TYPE63_REG          = 32'h100;
localparam JUMP_TYPE64_REG          = 32'h104;
localparam JUMP_TYPE65_REG          = 32'h108;
localparam JUMP_TYPE66_REG          = 32'h10c;
localparam JUMP_TYPE67_REG          = 32'h110;
localparam JUMP_TYPE68_REG          = 32'h114;
localparam JUMP_TYPE69_REG          = 32'h118;
localparam JUMP_TYPE70_REG          = 32'h11c;
localparam JUMP_TYPE71_REG          = 32'h120;
localparam JUMP_TYPE72_REG          = 32'h124;
localparam JUMP_TYPE73_REG          = 32'h128;
localparam JUMP_TYPE74_REG          = 32'h12c;
localparam JUMP_TYPE75_REG          = 32'h130;
localparam JUMP_TYPE76_REG          = 32'h134;
localparam JUMP_TYPE77_REG          = 32'h138;
localparam JUMP_TYPE78_REG          = 32'h13c;
localparam JUMP_TYPE79_REG          = 32'h140;
localparam JUMP_TYPE80_REG          = 32'h144;
localparam JUMP_TYPE81_REG          = 32'h148;
localparam JUMP_TYPE82_REG          = 32'h14c;
localparam JUMP_TYPE83_REG          = 32'h150;
localparam JUMP_TYPE84_REG          = 32'h154;
localparam JUMP_TYPE85_REG          = 32'h158;
localparam JUMP_TYPE86_REG          = 32'h15c;
localparam JUMP_TYPE87_REG          = 32'h160;
localparam JUMP_TYPE88_REG          = 32'h164;
localparam JUMP_TYPE89_REG          = 32'h168;
localparam JUMP_TYPE90_REG          = 32'h16c;
localparam JUMP_TYPE91_REG          = 32'h170;
localparam JUMP_TYPE92_REG          = 32'h174;
localparam JUMP_TYPE93_REG          = 32'h178;
localparam JUMP_TYPE94_REG          = 32'h17c;
localparam JUMP_TYPE95_REG          = 32'h180;
localparam JUMP_TYPE96_REG          = 32'h184;
localparam JUMP_TYPE97_REG          = 32'h188;
localparam JUMP_TYPE98_REG          = 32'h18c;
localparam JUMP_TYPE99_REG          = 32'h190;
localparam JUMP_TYPE100_REG         = 32'h194;
localparam JUMP_TYPE101_REG         = 32'h198;
localparam JUMP_TYPE102_REG         = 32'h19c;
localparam JUMP_TYPE103_REG         = 32'h1a0;
localparam JUMP_TYPE104_REG         = 32'h1a4;
localparam JUMP_TYPE105_REG         = 32'h1a8;
localparam JUMP_TYPE106_REG         = 32'h1ac;
localparam JUMP_TYPE107_REG         = 32'h1b0;
localparam JUMP_TYPE108_REG         = 32'h1b4;
localparam JUMP_TYPE109_REG         = 32'h1b8;
localparam JUMP_TYPE110_REG         = 32'h1bc;
localparam JUMP_TYPE111_REG         = 32'h1c0;
localparam JUMP_TYPE112_REG         = 32'h1c4;
localparam JUMP_TYPE113_REG         = 32'h1c8;
localparam JUMP_TYPE114_REG         = 32'h1cc;
localparam JUMP_TYPE115_REG         = 32'h1d0;
localparam JUMP_TYPE116_REG         = 32'h1d4;
localparam JUMP_TYPE117_REG         = 32'h1d8;
localparam JUMP_TYPE118_REG         = 32'h1dc;
localparam JUMP_TYPE119_REG         = 32'h1e0;
localparam JUMP_TYPE120_REG         = 32'h1e4;
localparam JUMP_TYPE121_REG         = 32'h1e8;
localparam JUMP_TYPE122_REG         = 32'h1ec;
localparam JUMP_TYPE123_REG         = 32'h1f0;
localparam JUMP_TYPE124_REG         = 32'h1f4;
localparam JUMP_TYPE125_REG         = 32'h1f8;
localparam JUMP_TYPE126_REG         = 32'h1fc;
localparam JUMP_TYPE127_REG         = 32'h200;
localparam JUMP_TYPE128_REG         = 32'h204;
localparam JUMP_TYPE129_REG         = 32'h208;
localparam JUMP_TYPE130_REG         = 32'h20c;
localparam JUMP_TYPE131_REG         = 32'h210;
localparam JUMP_TYPE132_REG         = 32'h214;
localparam JUMP_TYPE133_REG         = 32'h218;
localparam JUMP_TYPE134_REG         = 32'h21c;
localparam JUMP_TYPE135_REG         = 32'h220;
localparam JUMP_TYPE136_REG         = 32'h224;
localparam JUMP_TYPE137_REG         = 32'h228;
localparam JUMP_TYPE138_REG         = 32'h22c;
localparam JUMP_TYPE139_REG         = 32'h230;
localparam JUMP_TYPE140_REG         = 32'h234;
localparam JUMP_TYPE141_REG         = 32'h238;
localparam JUMP_TYPE142_REG         = 32'h23c;
localparam JUMP_TYPE143_REG         = 32'h240;
localparam JUMP_TYPE144_REG         = 32'h244;
localparam JUMP_TYPE145_REG         = 32'h248;
localparam JUMP_TYPE146_REG         = 32'h24c;
localparam JUMP_TYPE147_REG         = 32'h250;
localparam JUMP_TYPE148_REG         = 32'h254;
localparam JUMP_TYPE149_REG         = 32'h258;
localparam JUMP_TYPE150_REG         = 32'h25c;
localparam JUMP_TYPE151_REG         = 32'h260;
localparam JUMP_TYPE152_REG         = 32'h264;
localparam JUMP_TYPE153_REG         = 32'h268;
localparam JUMP_TYPE154_REG         = 32'h26c;
localparam JUMP_TYPE155_REG         = 32'h270;
localparam JUMP_TYPE156_REG         = 32'h274;
localparam JUMP_TYPE157_REG         = 32'h278;
localparam JUMP_TYPE158_REG         = 32'h27c;
localparam JUMP_TYPE159_REG         = 32'h280;
localparam JUMP_TYPE160_REG         = 32'h284;
localparam JUMP_TYPE161_REG         = 32'h288;
localparam JUMP_TYPE162_REG         = 32'h28c;
localparam JUMP_TYPE163_REG         = 32'h290;
localparam JUMP_TYPE164_REG         = 32'h294;
localparam JUMP_TYPE165_REG         = 32'h298;
localparam JUMP_TYPE166_REG         = 32'h29c;
localparam JUMP_TYPE167_REG         = 32'h2a0;
localparam JUMP_TYPE168_REG         = 32'h2a4;
localparam JUMP_TYPE169_REG         = 32'h2a8;
localparam JUMP_TYPE170_REG         = 32'h2ac;
localparam JUMP_TYPE171_REG         = 32'h2b0;
localparam JUMP_TYPE172_REG         = 32'h2b4;
localparam JUMP_TYPE173_REG         = 32'h2b8;
localparam JUMP_TYPE174_REG         = 32'h2bc;
localparam JUMP_TYPE175_REG         = 32'h2c0;
localparam JUMP_TYPE176_REG         = 32'h2c4;
localparam JUMP_TYPE177_REG         = 32'h2c8;
localparam JUMP_TYPE178_REG         = 32'h2cc;
localparam JUMP_TYPE179_REG         = 32'h2d0;
localparam JUMP_TYPE180_REG         = 32'h2d4;
localparam JUMP_TYPE181_REG         = 32'h2d8;
localparam JUMP_TYPE182_REG         = 32'h2dc;
localparam JUMP_TYPE183_REG         = 32'h2e0;
localparam JUMP_TYPE184_REG         = 32'h2e4;
localparam JUMP_TYPE185_REG         = 32'h2e8;
localparam JUMP_TYPE186_REG         = 32'h2ec;
localparam JUMP_TYPE187_REG         = 32'h2f0;
localparam JUMP_TYPE188_REG         = 32'h2f4;
localparam JUMP_TYPE189_REG         = 32'h2f8;
localparam JUMP_TYPE190_REG         = 32'h2fc;
localparam JUMP_TYPE191_REG         = 32'h300;
localparam JUMP_TYPE192_REG         = 32'h304;
localparam JUMP_TYPE193_REG         = 32'h308;
localparam JUMP_TYPE194_REG         = 32'h30c;
localparam JUMP_TYPE195_REG         = 32'h310;
localparam JUMP_TYPE196_REG         = 32'h314;
localparam JUMP_TYPE197_REG         = 32'h318;
localparam JUMP_TYPE198_REG         = 32'h31c;
localparam JUMP_TYPE199_REG         = 32'h320;
localparam JUMP_TYPE200_REG         = 32'h324;
localparam JUMP_TYPE201_REG         = 32'h328;
localparam JUMP_TYPE202_REG         = 32'h32c;
localparam JUMP_TYPE203_REG         = 32'h330;
localparam JUMP_TYPE204_REG         = 32'h334;
localparam JUMP_TYPE205_REG         = 32'h338;
localparam JUMP_TYPE206_REG         = 32'h33c;
localparam JUMP_TYPE207_REG         = 32'h340;
localparam JUMP_TYPE208_REG         = 32'h344;
localparam JUMP_TYPE209_REG         = 32'h348;
localparam JUMP_TYPE210_REG         = 32'h34c;
localparam JUMP_TYPE211_REG         = 32'h350;
localparam JUMP_TYPE212_REG         = 32'h354;
localparam JUMP_TYPE213_REG         = 32'h358;
localparam JUMP_TYPE214_REG         = 32'h35c;
localparam JUMP_TYPE215_REG         = 32'h360;
localparam JUMP_TYPE216_REG         = 32'h364;
localparam JUMP_TYPE217_REG         = 32'h368;
localparam JUMP_TYPE218_REG         = 32'h36c;
localparam JUMP_TYPE219_REG         = 32'h370;
localparam JUMP_TYPE220_REG         = 32'h374;
localparam JUMP_TYPE221_REG         = 32'h378;
localparam JUMP_TYPE222_REG         = 32'h37c;
localparam JUMP_TYPE223_REG         = 32'h380;
localparam JUMP_TYPE224_REG         = 32'h384;
localparam JUMP_TYPE225_REG         = 32'h388;
localparam JUMP_TYPE226_REG         = 32'h38c;
localparam JUMP_TYPE227_REG         = 32'h390;
localparam JUMP_TYPE228_REG         = 32'h394;
localparam JUMP_TYPE229_REG         = 32'h398;
localparam JUMP_TYPE230_REG         = 32'h39c;
localparam JUMP_TYPE231_REG         = 32'h3a0;
localparam JUMP_TYPE232_REG         = 32'h3a4;
localparam JUMP_TYPE233_REG         = 32'h3a8;
localparam JUMP_TYPE234_REG         = 32'h3ac;
localparam JUMP_TYPE235_REG         = 32'h3b0;
localparam JUMP_TYPE236_REG         = 32'h3b4;
localparam JUMP_TYPE237_REG         = 32'h3b8;
localparam JUMP_TYPE238_REG         = 32'h3bc;
localparam JUMP_TYPE239_REG         = 32'h3c0;
localparam JUMP_TYPE240_REG         = 32'h3c4;
localparam JUMP_TYPE241_REG         = 32'h3c8;
localparam JUMP_TYPE242_REG         = 32'h3cc;
localparam JUMP_TYPE243_REG         = 32'h3d0;
localparam JUMP_TYPE244_REG         = 32'h3d4;
localparam JUMP_TYPE245_REG         = 32'h3d8;
localparam JUMP_TYPE246_REG         = 32'h3dc;
localparam JUMP_TYPE247_REG         = 32'h3e0;
localparam JUMP_TYPE248_REG         = 32'h3e4;
localparam JUMP_TYPE249_REG         = 32'h3e8;
localparam JUMP_TYPE250_REG         = 32'h3ec;
localparam JUMP_TYPE251_REG         = 32'h3f0;
localparam JUMP_TYPE252_REG         = 32'h3f4;
localparam JUMP_TYPE253_REG         = 32'h3f8;
localparam JUMP_TYPE254_REG         = 32'h3fc;
localparam JUMP_TYPE255_REG         = 32'h400;
localparam JUMP_TYPE256_REG         = 32'h404;
localparam JUMP_TYPE257_REG         = 32'h408;
localparam JUMP_TYPE258_REG         = 32'h40c;
localparam JUMP_TYPE259_REG         = 32'h410;
localparam JUMP_TYPE260_REG         = 32'h414;
localparam JUMP_TYPE261_REG         = 32'h418;
localparam JUMP_TYPE262_REG         = 32'h41c;
localparam JUMP_TYPE263_REG         = 32'h420;
localparam JUMP_TYPE264_REG         = 32'h424;
localparam JUMP_TYPE265_REG         = 32'h428;
localparam JUMP_TYPE266_REG         = 32'h42c;
localparam JUMP_TYPE267_REG         = 32'h430;
localparam JUMP_TYPE268_REG         = 32'h434;
localparam JUMP_TYPE269_REG         = 32'h438;
localparam JUMP_TYPE270_REG         = 32'h43c;
localparam JUMP_TYPE271_REG         = 32'h440;
localparam JUMP_TYPE272_REG         = 32'h444;
localparam JUMP_TYPE273_REG         = 32'h448;
localparam JUMP_TYPE274_REG         = 32'h44c;
localparam JUMP_TYPE275_REG         = 32'h450;
localparam JUMP_TYPE276_REG         = 32'h454;
localparam JUMP_TYPE277_REG         = 32'h458;
localparam JUMP_TYPE278_REG         = 32'h45c;
localparam JUMP_TYPE279_REG         = 32'h460;
localparam JUMP_TYPE280_REG         = 32'h464;
localparam JUMP_TYPE281_REG         = 32'h468;
localparam JUMP_TYPE282_REG         = 32'h46c;
localparam JUMP_TYPE283_REG         = 32'h470;
localparam JUMP_TYPE284_REG         = 32'h474;
localparam JUMP_TYPE285_REG         = 32'h478;
localparam JUMP_TYPE286_REG         = 32'h47c;
localparam JUMP_TYPE287_REG         = 32'h480;
localparam JUMP_TYPE288_REG         = 32'h484;
localparam JUMP_TYPE289_REG         = 32'h488;
localparam JUMP_TYPE290_REG         = 32'h48c;
localparam JUMP_TYPE291_REG         = 32'h490;
localparam JUMP_TYPE292_REG         = 32'h494;
localparam JUMP_TYPE293_REG         = 32'h498;
localparam JUMP_TYPE294_REG         = 32'h49c;
localparam JUMP_TYPE295_REG         = 32'h4a0;
localparam JUMP_TYPE296_REG         = 32'h4a4;
localparam JUMP_TYPE297_REG         = 32'h4a8;
localparam JUMP_TYPE298_REG         = 32'h4ac;
localparam JUMP_TYPE299_REG         = 32'h4b0;
localparam JUMP_TYPE300_REG         = 32'h4b4;
localparam JUMP_TYPE301_REG         = 32'h4b8;
localparam JUMP_TYPE302_REG         = 32'h4bc;
localparam JUMP_TYPE303_REG         = 32'h4c0;
localparam JUMP_TYPE304_REG         = 32'h4c4;
localparam JUMP_TYPE305_REG         = 32'h4c8;
localparam JUMP_TYPE306_REG         = 32'h4cc;
localparam JUMP_TYPE307_REG         = 32'h4d0;
localparam JUMP_TYPE308_REG         = 32'h4d4;
localparam JUMP_TYPE309_REG         = 32'h4d8;
localparam JUMP_TYPE310_REG         = 32'h4dc;
localparam JUMP_TYPE311_REG         = 32'h4e0;
localparam JUMP_TYPE312_REG         = 32'h4e4;
localparam JUMP_TYPE313_REG         = 32'h4e8;
localparam JUMP_TYPE314_REG         = 32'h4ec;
localparam JUMP_TYPE315_REG         = 32'h4f0;
localparam JUMP_TYPE316_REG         = 32'h4f4;
localparam JUMP_TYPE317_REG         = 32'h4f8;
localparam JUMP_TYPE318_REG         = 32'h4fc;
localparam JUMP_TYPE319_REG         = 32'h500;
localparam JUMP_TYPE320_REG         = 32'h504;
localparam JUMP_TYPE321_REG         = 32'h508;
localparam JUMP_TYPE322_REG         = 32'h50c;
localparam JUMP_TYPE323_REG         = 32'h510;
localparam JUMP_TYPE324_REG         = 32'h514;
localparam JUMP_TYPE325_REG         = 32'h518;
localparam JUMP_TYPE326_REG         = 32'h51c;
localparam JUMP_TYPE327_REG         = 32'h520;
localparam JUMP_TYPE328_REG         = 32'h524;
localparam JUMP_TYPE329_REG         = 32'h528;
localparam JUMP_TYPE330_REG         = 32'h52c;
localparam JUMP_TYPE331_REG         = 32'h530;
localparam JUMP_TYPE332_REG         = 32'h534;
localparam JUMP_TYPE333_REG         = 32'h538;
localparam JUMP_TYPE334_REG         = 32'h53c;
localparam JUMP_TYPE335_REG         = 32'h540;
localparam JUMP_TYPE336_REG         = 32'h544;
localparam JUMP_TYPE337_REG         = 32'h548;
localparam JUMP_TYPE338_REG         = 32'h54c;
localparam JUMP_TYPE339_REG         = 32'h550;
localparam JUMP_TYPE340_REG         = 32'h554;
localparam JUMP_TYPE341_REG         = 32'h558;
localparam JUMP_TYPE342_REG         = 32'h55c;
localparam JUMP_TYPE343_REG         = 32'h560;
localparam JUMP_TYPE344_REG         = 32'h564;
localparam JUMP_TYPE345_REG         = 32'h568;
localparam JUMP_TYPE346_REG         = 32'h56c;
localparam JUMP_TYPE347_REG         = 32'h570;
localparam JUMP_TYPE348_REG         = 32'h574;
localparam JUMP_TYPE349_REG         = 32'h578;
localparam JUMP_TYPE350_REG         = 32'h57c;
localparam JUMP_TYPE351_REG         = 32'h580;
localparam JUMP_TYPE352_REG         = 32'h584;
localparam JUMP_TYPE353_REG         = 32'h588;
localparam JUMP_TYPE354_REG         = 32'h58c;
localparam JUMP_TYPE355_REG         = 32'h590;
localparam JUMP_TYPE356_REG         = 32'h594;
localparam JUMP_TYPE357_REG         = 32'h598;
localparam JUMP_TYPE358_REG         = 32'h59c;
localparam JUMP_TYPE359_REG         = 32'h5a0;
localparam JUMP_TYPE360_REG         = 32'h5a4;
localparam JUMP_TYPE361_REG         = 32'h5a8;
localparam JUMP_TYPE362_REG         = 32'h5ac;
localparam JUMP_TYPE363_REG         = 32'h5b0;
localparam JUMP_TYPE364_REG         = 32'h5b4;
localparam JUMP_TYPE365_REG         = 32'h5b8;
localparam JUMP_TYPE366_REG         = 32'h5bc;
localparam JUMP_TYPE367_REG         = 32'h5c0;
localparam JUMP_TYPE368_REG         = 32'h5c4;
localparam JUMP_TYPE369_REG         = 32'h5c8;
localparam JUMP_TYPE370_REG         = 32'h5cc;
localparam JUMP_TYPE371_REG         = 32'h5d0;
localparam JUMP_TYPE372_REG         = 32'h5d4;
localparam JUMP_TYPE373_REG         = 32'h5d8;
localparam JUMP_TYPE374_REG         = 32'h5dc;
localparam JUMP_TYPE375_REG         = 32'h5e0;
localparam JUMP_TYPE376_REG         = 32'h5e4;
localparam JUMP_TYPE377_REG         = 32'h5e8;
localparam JUMP_TYPE378_REG         = 32'h5ec;
localparam JUMP_TYPE379_REG         = 32'h5f0;
localparam JUMP_TYPE380_REG         = 32'h5f4;
localparam JUMP_TYPE381_REG         = 32'h5f8;
localparam JUMP_TYPE382_REG         = 32'h5fc;
localparam JUMP_TYPE383_REG         = 32'h600;
localparam JUMP_TYPE384_REG         = 32'h604;
localparam JUMP_TYPE385_REG         = 32'h608;
localparam JUMP_TYPE386_REG         = 32'h60c;
localparam JUMP_TYPE387_REG         = 32'h610;
localparam JUMP_TYPE388_REG         = 32'h614;
localparam JUMP_TYPE389_REG         = 32'h618;
localparam JUMP_TYPE390_REG         = 32'h61c;
localparam JUMP_TYPE391_REG         = 32'h620;
localparam JUMP_TYPE392_REG         = 32'h624;
localparam JUMP_TYPE393_REG         = 32'h628;
localparam JUMP_TYPE394_REG         = 32'h62c;
localparam JUMP_TYPE395_REG         = 32'h630;
localparam JUMP_TYPE396_REG         = 32'h634;
localparam JUMP_TYPE397_REG         = 32'h638;
localparam JUMP_TYPE398_REG         = 32'h63c;
localparam JUMP_TYPE399_REG         = 32'h640;
localparam JUMP_TYPE400_REG         = 32'h644;
localparam JUMP_TYPE401_REG         = 32'h648;
localparam JUMP_TYPE402_REG         = 32'h64c;
localparam JUMP_TYPE403_REG         = 32'h650;
localparam JUMP_TYPE404_REG         = 32'h654;
localparam JUMP_TYPE405_REG         = 32'h658;
localparam JUMP_TYPE406_REG         = 32'h65c;
localparam JUMP_TYPE407_REG         = 32'h660;
localparam JUMP_TYPE408_REG         = 32'h664;
localparam JUMP_TYPE409_REG         = 32'h668;
localparam JUMP_TYPE410_REG         = 32'h66c;
localparam JUMP_TYPE411_REG         = 32'h670;
localparam JUMP_TYPE412_REG         = 32'h674;
localparam JUMP_TYPE413_REG         = 32'h678;
localparam JUMP_TYPE414_REG         = 32'h67c;
localparam JUMP_TYPE415_REG         = 32'h680;
localparam JUMP_TYPE416_REG         = 32'h684;
localparam JUMP_TYPE417_REG         = 32'h688;
localparam JUMP_TYPE418_REG         = 32'h68c;
localparam JUMP_TYPE419_REG         = 32'h690;
localparam JUMP_TYPE420_REG         = 32'h694;
localparam JUMP_TYPE421_REG         = 32'h698;
localparam JUMP_TYPE422_REG         = 32'h69c;
localparam JUMP_TYPE423_REG         = 32'h6a0;
localparam JUMP_TYPE424_REG         = 32'h6a4;
localparam JUMP_TYPE425_REG         = 32'h6a8;
localparam JUMP_TYPE426_REG         = 32'h6ac;
localparam JUMP_TYPE427_REG         = 32'h6b0;
localparam JUMP_TYPE428_REG         = 32'h6b4;
localparam JUMP_TYPE429_REG         = 32'h6b8;
localparam JUMP_TYPE430_REG         = 32'h6bc;
localparam JUMP_TYPE431_REG         = 32'h6c0;
localparam JUMP_TYPE432_REG         = 32'h6c4;
localparam JUMP_TYPE433_REG         = 32'h6c8;
localparam JUMP_TYPE434_REG         = 32'h6cc;
localparam JUMP_TYPE435_REG         = 32'h6d0;
localparam JUMP_TYPE436_REG         = 32'h6d4;
localparam JUMP_TYPE437_REG         = 32'h6d8;
localparam JUMP_TYPE438_REG         = 32'h6dc;
localparam JUMP_TYPE439_REG         = 32'h6e0;
localparam JUMP_TYPE440_REG         = 32'h6e4;
localparam JUMP_TYPE441_REG         = 32'h6e8;
localparam JUMP_TYPE442_REG         = 32'h6ec;
localparam JUMP_TYPE443_REG         = 32'h6f0;
localparam JUMP_TYPE444_REG         = 32'h6f4;
localparam JUMP_TYPE445_REG         = 32'h6f8;
localparam JUMP_TYPE446_REG         = 32'h6fc;
localparam JUMP_TYPE447_REG         = 32'h700;
localparam JUMP_TYPE448_REG         = 32'h704;
localparam JUMP_TYPE449_REG         = 32'h708;
localparam JUMP_TYPE450_REG         = 32'h70c;
localparam JUMP_TYPE451_REG         = 32'h710;
localparam JUMP_TYPE452_REG         = 32'h714;
localparam JUMP_TYPE453_REG         = 32'h718;
localparam JUMP_TYPE454_REG         = 32'h71c;
localparam JUMP_TYPE455_REG         = 32'h720;
localparam JUMP_TYPE456_REG         = 32'h724;
localparam JUMP_TYPE457_REG         = 32'h728;
localparam JUMP_TYPE458_REG         = 32'h72c;
localparam JUMP_TYPE459_REG         = 32'h730;
localparam JUMP_TYPE460_REG         = 32'h734;
localparam JUMP_TYPE461_REG         = 32'h738;
localparam JUMP_TYPE462_REG         = 32'h73c;
localparam JUMP_TYPE463_REG         = 32'h740;
localparam JUMP_TYPE464_REG         = 32'h744;
localparam JUMP_TYPE465_REG         = 32'h748;
localparam JUMP_TYPE466_REG         = 32'h74c;
localparam JUMP_TYPE467_REG         = 32'h750;
localparam JUMP_TYPE468_REG         = 32'h754;
localparam JUMP_TYPE469_REG         = 32'h758;
localparam JUMP_TYPE470_REG         = 32'h75c;
localparam JUMP_TYPE471_REG         = 32'h760;
localparam JUMP_TYPE472_REG         = 32'h764;
localparam JUMP_TYPE473_REG         = 32'h768;
localparam JUMP_TYPE474_REG         = 32'h76c;
localparam JUMP_TYPE475_REG         = 32'h770;
localparam JUMP_TYPE476_REG         = 32'h774;
localparam JUMP_TYPE477_REG         = 32'h778;
localparam JUMP_TYPE478_REG         = 32'h77c;
localparam JUMP_TYPE479_REG         = 32'h780;
localparam JUMP_TYPE480_REG         = 32'h784;
localparam JUMP_TYPE481_REG         = 32'h788;
localparam JUMP_TYPE482_REG         = 32'h78c;
localparam JUMP_TYPE483_REG         = 32'h790;
localparam JUMP_TYPE484_REG         = 32'h794;
localparam JUMP_TYPE485_REG         = 32'h798;
localparam JUMP_TYPE486_REG         = 32'h79c;
localparam JUMP_TYPE487_REG         = 32'h7a0;
localparam JUMP_TYPE488_REG         = 32'h7a4;
localparam JUMP_TYPE489_REG         = 32'h7a8;
localparam JUMP_TYPE490_REG         = 32'h7ac;
localparam JUMP_TYPE491_REG         = 32'h7b0;
localparam JUMP_TYPE492_REG         = 32'h7b4;
localparam JUMP_TYPE493_REG         = 32'h7b8;
localparam JUMP_TYPE494_REG         = 32'h7bc;
localparam JUMP_TYPE495_REG         = 32'h7c0;
localparam JUMP_TYPE496_REG         = 32'h7c4;
localparam JUMP_TYPE497_REG         = 32'h7c8;
localparam JUMP_TYPE498_REG         = 32'h7cc;
localparam JUMP_TYPE499_REG         = 32'h7d0;
localparam JUMP_TYPE500_REG         = 32'h7d4;
localparam JUMP_TYPE501_REG         = 32'h7d8;
localparam JUMP_TYPE502_REG         = 32'h7dc;
localparam JUMP_TYPE503_REG         = 32'h7e0;
localparam JUMP_TYPE504_REG         = 32'h7e4;
localparam JUMP_TYPE505_REG         = 32'h7e8;
localparam JUMP_TYPE506_REG         = 32'h7ec;
localparam JUMP_TYPE507_REG         = 32'h7f0;
localparam JUMP_TYPE508_REG         = 32'h7f4;
localparam JUMP_TYPE509_REG         = 32'h7f8;
localparam JUMP_TYPE510_REG         = 32'h7fc;
localparam JUMP_TYPE511_REG         = 32'h800;

//----------------------------local wire/reg declaration------------------------------------------
wire [32-1:0] common_para_reg             ;
wire [32-1:0] jump_type0_reg              ;
wire [32-1:0] jump_type1_reg              ;
wire [32-1:0] jump_type2_reg              ;
wire [32-1:0] jump_type3_reg              ;
wire [32-1:0] jump_type4_reg              ;
wire [32-1:0] jump_type5_reg              ;
wire [32-1:0] jump_type6_reg              ;
wire [32-1:0] jump_type7_reg              ;
wire [32-1:0] jump_type8_reg              ;
wire [32-1:0] jump_type9_reg              ;
wire [32-1:0] jump_type10_reg             ;
wire [32-1:0] jump_type11_reg             ;
wire [32-1:0] jump_type12_reg             ;
wire [32-1:0] jump_type13_reg             ;
wire [32-1:0] jump_type14_reg             ;
wire [32-1:0] jump_type15_reg             ;
wire [32-1:0] jump_type16_reg             ;
wire [32-1:0] jump_type17_reg             ;
wire [32-1:0] jump_type18_reg             ;
wire [32-1:0] jump_type19_reg             ;
wire [32-1:0] jump_type20_reg             ;
wire [32-1:0] jump_type21_reg             ;
wire [32-1:0] jump_type22_reg             ;
wire [32-1:0] jump_type23_reg             ;
wire [32-1:0] jump_type24_reg             ;
wire [32-1:0] jump_type25_reg             ;
wire [32-1:0] jump_type26_reg             ;
wire [32-1:0] jump_type27_reg             ;
wire [32-1:0] jump_type28_reg             ;
wire [32-1:0] jump_type29_reg             ;
wire [32-1:0] jump_type30_reg             ;
wire [32-1:0] jump_type31_reg             ;
wire [32-1:0] jump_type32_reg             ;
wire [32-1:0] jump_type33_reg             ;
wire [32-1:0] jump_type34_reg             ;
wire [32-1:0] jump_type35_reg             ;
wire [32-1:0] jump_type36_reg             ;
wire [32-1:0] jump_type37_reg             ;
wire [32-1:0] jump_type38_reg             ;
wire [32-1:0] jump_type39_reg             ;
wire [32-1:0] jump_type40_reg             ;
wire [32-1:0] jump_type41_reg             ;
wire [32-1:0] jump_type42_reg             ;
wire [32-1:0] jump_type43_reg             ;
wire [32-1:0] jump_type44_reg             ;
wire [32-1:0] jump_type45_reg             ;
wire [32-1:0] jump_type46_reg             ;
wire [32-1:0] jump_type47_reg             ;
wire [32-1:0] jump_type48_reg             ;
wire [32-1:0] jump_type49_reg             ;
wire [32-1:0] jump_type50_reg             ;
wire [32-1:0] jump_type51_reg             ;
wire [32-1:0] jump_type52_reg             ;
wire [32-1:0] jump_type53_reg             ;
wire [32-1:0] jump_type54_reg             ;
wire [32-1:0] jump_type55_reg             ;
wire [32-1:0] jump_type56_reg             ;
wire [32-1:0] jump_type57_reg             ;
wire [32-1:0] jump_type58_reg             ;
wire [32-1:0] jump_type59_reg             ;
wire [32-1:0] jump_type60_reg             ;
wire [32-1:0] jump_type61_reg             ;
wire [32-1:0] jump_type62_reg             ;
wire [32-1:0] jump_type63_reg             ;
wire [32-1:0] jump_type64_reg             ;
wire [32-1:0] jump_type65_reg             ;
wire [32-1:0] jump_type66_reg             ;
wire [32-1:0] jump_type67_reg             ;
wire [32-1:0] jump_type68_reg             ;
wire [32-1:0] jump_type69_reg             ;
wire [32-1:0] jump_type70_reg             ;
wire [32-1:0] jump_type71_reg             ;
wire [32-1:0] jump_type72_reg             ;
wire [32-1:0] jump_type73_reg             ;
wire [32-1:0] jump_type74_reg             ;
wire [32-1:0] jump_type75_reg             ;
wire [32-1:0] jump_type76_reg             ;
wire [32-1:0] jump_type77_reg             ;
wire [32-1:0] jump_type78_reg             ;
wire [32-1:0] jump_type79_reg             ;
wire [32-1:0] jump_type80_reg             ;
wire [32-1:0] jump_type81_reg             ;
wire [32-1:0] jump_type82_reg             ;
wire [32-1:0] jump_type83_reg             ;
wire [32-1:0] jump_type84_reg             ;
wire [32-1:0] jump_type85_reg             ;
wire [32-1:0] jump_type86_reg             ;
wire [32-1:0] jump_type87_reg             ;
wire [32-1:0] jump_type88_reg             ;
wire [32-1:0] jump_type89_reg             ;
wire [32-1:0] jump_type90_reg             ;
wire [32-1:0] jump_type91_reg             ;
wire [32-1:0] jump_type92_reg             ;
wire [32-1:0] jump_type93_reg             ;
wire [32-1:0] jump_type94_reg             ;
wire [32-1:0] jump_type95_reg             ;
wire [32-1:0] jump_type96_reg             ;
wire [32-1:0] jump_type97_reg             ;
wire [32-1:0] jump_type98_reg             ;
wire [32-1:0] jump_type99_reg             ;
wire [32-1:0] jump_type100_reg            ;
wire [32-1:0] jump_type101_reg            ;
wire [32-1:0] jump_type102_reg            ;
wire [32-1:0] jump_type103_reg            ;
wire [32-1:0] jump_type104_reg            ;
wire [32-1:0] jump_type105_reg            ;
wire [32-1:0] jump_type106_reg            ;
wire [32-1:0] jump_type107_reg            ;
wire [32-1:0] jump_type108_reg            ;
wire [32-1:0] jump_type109_reg            ;
wire [32-1:0] jump_type110_reg            ;
wire [32-1:0] jump_type111_reg            ;
wire [32-1:0] jump_type112_reg            ;
wire [32-1:0] jump_type113_reg            ;
wire [32-1:0] jump_type114_reg            ;
wire [32-1:0] jump_type115_reg            ;
wire [32-1:0] jump_type116_reg            ;
wire [32-1:0] jump_type117_reg            ;
wire [32-1:0] jump_type118_reg            ;
wire [32-1:0] jump_type119_reg            ;
wire [32-1:0] jump_type120_reg            ;
wire [32-1:0] jump_type121_reg            ;
wire [32-1:0] jump_type122_reg            ;
wire [32-1:0] jump_type123_reg            ;
wire [32-1:0] jump_type124_reg            ;
wire [32-1:0] jump_type125_reg            ;
wire [32-1:0] jump_type126_reg            ;
wire [32-1:0] jump_type127_reg            ;
wire [32-1:0] jump_type128_reg            ;
wire [32-1:0] jump_type129_reg            ;
wire [32-1:0] jump_type130_reg            ;
wire [32-1:0] jump_type131_reg            ;
wire [32-1:0] jump_type132_reg            ;
wire [32-1:0] jump_type133_reg            ;
wire [32-1:0] jump_type134_reg            ;
wire [32-1:0] jump_type135_reg            ;
wire [32-1:0] jump_type136_reg            ;
wire [32-1:0] jump_type137_reg            ;
wire [32-1:0] jump_type138_reg            ;
wire [32-1:0] jump_type139_reg            ;
wire [32-1:0] jump_type140_reg            ;
wire [32-1:0] jump_type141_reg            ;
wire [32-1:0] jump_type142_reg            ;
wire [32-1:0] jump_type143_reg            ;
wire [32-1:0] jump_type144_reg            ;
wire [32-1:0] jump_type145_reg            ;
wire [32-1:0] jump_type146_reg            ;
wire [32-1:0] jump_type147_reg            ;
wire [32-1:0] jump_type148_reg            ;
wire [32-1:0] jump_type149_reg            ;
wire [32-1:0] jump_type150_reg            ;
wire [32-1:0] jump_type151_reg            ;
wire [32-1:0] jump_type152_reg            ;
wire [32-1:0] jump_type153_reg            ;
wire [32-1:0] jump_type154_reg            ;
wire [32-1:0] jump_type155_reg            ;
wire [32-1:0] jump_type156_reg            ;
wire [32-1:0] jump_type157_reg            ;
wire [32-1:0] jump_type158_reg            ;
wire [32-1:0] jump_type159_reg            ;
wire [32-1:0] jump_type160_reg            ;
wire [32-1:0] jump_type161_reg            ;
wire [32-1:0] jump_type162_reg            ;
wire [32-1:0] jump_type163_reg            ;
wire [32-1:0] jump_type164_reg            ;
wire [32-1:0] jump_type165_reg            ;
wire [32-1:0] jump_type166_reg            ;
wire [32-1:0] jump_type167_reg            ;
wire [32-1:0] jump_type168_reg            ;
wire [32-1:0] jump_type169_reg            ;
wire [32-1:0] jump_type170_reg            ;
wire [32-1:0] jump_type171_reg            ;
wire [32-1:0] jump_type172_reg            ;
wire [32-1:0] jump_type173_reg            ;
wire [32-1:0] jump_type174_reg            ;
wire [32-1:0] jump_type175_reg            ;
wire [32-1:0] jump_type176_reg            ;
wire [32-1:0] jump_type177_reg            ;
wire [32-1:0] jump_type178_reg            ;
wire [32-1:0] jump_type179_reg            ;
wire [32-1:0] jump_type180_reg            ;
wire [32-1:0] jump_type181_reg            ;
wire [32-1:0] jump_type182_reg            ;
wire [32-1:0] jump_type183_reg            ;
wire [32-1:0] jump_type184_reg            ;
wire [32-1:0] jump_type185_reg            ;
wire [32-1:0] jump_type186_reg            ;
wire [32-1:0] jump_type187_reg            ;
wire [32-1:0] jump_type188_reg            ;
wire [32-1:0] jump_type189_reg            ;
wire [32-1:0] jump_type190_reg            ;
wire [32-1:0] jump_type191_reg            ;
wire [32-1:0] jump_type192_reg            ;
wire [32-1:0] jump_type193_reg            ;
wire [32-1:0] jump_type194_reg            ;
wire [32-1:0] jump_type195_reg            ;
wire [32-1:0] jump_type196_reg            ;
wire [32-1:0] jump_type197_reg            ;
wire [32-1:0] jump_type198_reg            ;
wire [32-1:0] jump_type199_reg            ;
wire [32-1:0] jump_type200_reg            ;
wire [32-1:0] jump_type201_reg            ;
wire [32-1:0] jump_type202_reg            ;
wire [32-1:0] jump_type203_reg            ;
wire [32-1:0] jump_type204_reg            ;
wire [32-1:0] jump_type205_reg            ;
wire [32-1:0] jump_type206_reg            ;
wire [32-1:0] jump_type207_reg            ;
wire [32-1:0] jump_type208_reg            ;
wire [32-1:0] jump_type209_reg            ;
wire [32-1:0] jump_type210_reg            ;
wire [32-1:0] jump_type211_reg            ;
wire [32-1:0] jump_type212_reg            ;
wire [32-1:0] jump_type213_reg            ;
wire [32-1:0] jump_type214_reg            ;
wire [32-1:0] jump_type215_reg            ;
wire [32-1:0] jump_type216_reg            ;
wire [32-1:0] jump_type217_reg            ;
wire [32-1:0] jump_type218_reg            ;
wire [32-1:0] jump_type219_reg            ;
wire [32-1:0] jump_type220_reg            ;
wire [32-1:0] jump_type221_reg            ;
wire [32-1:0] jump_type222_reg            ;
wire [32-1:0] jump_type223_reg            ;
wire [32-1:0] jump_type224_reg            ;
wire [32-1:0] jump_type225_reg            ;
wire [32-1:0] jump_type226_reg            ;
wire [32-1:0] jump_type227_reg            ;
wire [32-1:0] jump_type228_reg            ;
wire [32-1:0] jump_type229_reg            ;
wire [32-1:0] jump_type230_reg            ;
wire [32-1:0] jump_type231_reg            ;
wire [32-1:0] jump_type232_reg            ;
wire [32-1:0] jump_type233_reg            ;
wire [32-1:0] jump_type234_reg            ;
wire [32-1:0] jump_type235_reg            ;
wire [32-1:0] jump_type236_reg            ;
wire [32-1:0] jump_type237_reg            ;
wire [32-1:0] jump_type238_reg            ;
wire [32-1:0] jump_type239_reg            ;
wire [32-1:0] jump_type240_reg            ;
wire [32-1:0] jump_type241_reg            ;
wire [32-1:0] jump_type242_reg            ;
wire [32-1:0] jump_type243_reg            ;
wire [32-1:0] jump_type244_reg            ;
wire [32-1:0] jump_type245_reg            ;
wire [32-1:0] jump_type246_reg            ;
wire [32-1:0] jump_type247_reg            ;
wire [32-1:0] jump_type248_reg            ;
wire [32-1:0] jump_type249_reg            ;
wire [32-1:0] jump_type250_reg            ;
wire [32-1:0] jump_type251_reg            ;
wire [32-1:0] jump_type252_reg            ;
wire [32-1:0] jump_type253_reg            ;
wire [32-1:0] jump_type254_reg            ;
wire [32-1:0] jump_type255_reg            ;
wire [32-1:0] jump_type256_reg            ;
wire [32-1:0] jump_type257_reg            ;
wire [32-1:0] jump_type258_reg            ;
wire [32-1:0] jump_type259_reg            ;
wire [32-1:0] jump_type260_reg            ;
wire [32-1:0] jump_type261_reg            ;
wire [32-1:0] jump_type262_reg            ;
wire [32-1:0] jump_type263_reg            ;
wire [32-1:0] jump_type264_reg            ;
wire [32-1:0] jump_type265_reg            ;
wire [32-1:0] jump_type266_reg            ;
wire [32-1:0] jump_type267_reg            ;
wire [32-1:0] jump_type268_reg            ;
wire [32-1:0] jump_type269_reg            ;
wire [32-1:0] jump_type270_reg            ;
wire [32-1:0] jump_type271_reg            ;
wire [32-1:0] jump_type272_reg            ;
wire [32-1:0] jump_type273_reg            ;
wire [32-1:0] jump_type274_reg            ;
wire [32-1:0] jump_type275_reg            ;
wire [32-1:0] jump_type276_reg            ;
wire [32-1:0] jump_type277_reg            ;
wire [32-1:0] jump_type278_reg            ;
wire [32-1:0] jump_type279_reg            ;
wire [32-1:0] jump_type280_reg            ;
wire [32-1:0] jump_type281_reg            ;
wire [32-1:0] jump_type282_reg            ;
wire [32-1:0] jump_type283_reg            ;
wire [32-1:0] jump_type284_reg            ;
wire [32-1:0] jump_type285_reg            ;
wire [32-1:0] jump_type286_reg            ;
wire [32-1:0] jump_type287_reg            ;
wire [32-1:0] jump_type288_reg            ;
wire [32-1:0] jump_type289_reg            ;
wire [32-1:0] jump_type290_reg            ;
wire [32-1:0] jump_type291_reg            ;
wire [32-1:0] jump_type292_reg            ;
wire [32-1:0] jump_type293_reg            ;
wire [32-1:0] jump_type294_reg            ;
wire [32-1:0] jump_type295_reg            ;
wire [32-1:0] jump_type296_reg            ;
wire [32-1:0] jump_type297_reg            ;
wire [32-1:0] jump_type298_reg            ;
wire [32-1:0] jump_type299_reg            ;
wire [32-1:0] jump_type300_reg            ;
wire [32-1:0] jump_type301_reg            ;
wire [32-1:0] jump_type302_reg            ;
wire [32-1:0] jump_type303_reg            ;
wire [32-1:0] jump_type304_reg            ;
wire [32-1:0] jump_type305_reg            ;
wire [32-1:0] jump_type306_reg            ;
wire [32-1:0] jump_type307_reg            ;
wire [32-1:0] jump_type308_reg            ;
wire [32-1:0] jump_type309_reg            ;
wire [32-1:0] jump_type310_reg            ;
wire [32-1:0] jump_type311_reg            ;
wire [32-1:0] jump_type312_reg            ;
wire [32-1:0] jump_type313_reg            ;
wire [32-1:0] jump_type314_reg            ;
wire [32-1:0] jump_type315_reg            ;
wire [32-1:0] jump_type316_reg            ;
wire [32-1:0] jump_type317_reg            ;
wire [32-1:0] jump_type318_reg            ;
wire [32-1:0] jump_type319_reg            ;
wire [32-1:0] jump_type320_reg            ;
wire [32-1:0] jump_type321_reg            ;
wire [32-1:0] jump_type322_reg            ;
wire [32-1:0] jump_type323_reg            ;
wire [32-1:0] jump_type324_reg            ;
wire [32-1:0] jump_type325_reg            ;
wire [32-1:0] jump_type326_reg            ;
wire [32-1:0] jump_type327_reg            ;
wire [32-1:0] jump_type328_reg            ;
wire [32-1:0] jump_type329_reg            ;
wire [32-1:0] jump_type330_reg            ;
wire [32-1:0] jump_type331_reg            ;
wire [32-1:0] jump_type332_reg            ;
wire [32-1:0] jump_type333_reg            ;
wire [32-1:0] jump_type334_reg            ;
wire [32-1:0] jump_type335_reg            ;
wire [32-1:0] jump_type336_reg            ;
wire [32-1:0] jump_type337_reg            ;
wire [32-1:0] jump_type338_reg            ;
wire [32-1:0] jump_type339_reg            ;
wire [32-1:0] jump_type340_reg            ;
wire [32-1:0] jump_type341_reg            ;
wire [32-1:0] jump_type342_reg            ;
wire [32-1:0] jump_type343_reg            ;
wire [32-1:0] jump_type344_reg            ;
wire [32-1:0] jump_type345_reg            ;
wire [32-1:0] jump_type346_reg            ;
wire [32-1:0] jump_type347_reg            ;
wire [32-1:0] jump_type348_reg            ;
wire [32-1:0] jump_type349_reg            ;
wire [32-1:0] jump_type350_reg            ;
wire [32-1:0] jump_type351_reg            ;
wire [32-1:0] jump_type352_reg            ;
wire [32-1:0] jump_type353_reg            ;
wire [32-1:0] jump_type354_reg            ;
wire [32-1:0] jump_type355_reg            ;
wire [32-1:0] jump_type356_reg            ;
wire [32-1:0] jump_type357_reg            ;
wire [32-1:0] jump_type358_reg            ;
wire [32-1:0] jump_type359_reg            ;
wire [32-1:0] jump_type360_reg            ;
wire [32-1:0] jump_type361_reg            ;
wire [32-1:0] jump_type362_reg            ;
wire [32-1:0] jump_type363_reg            ;
wire [32-1:0] jump_type364_reg            ;
wire [32-1:0] jump_type365_reg            ;
wire [32-1:0] jump_type366_reg            ;
wire [32-1:0] jump_type367_reg            ;
wire [32-1:0] jump_type368_reg            ;
wire [32-1:0] jump_type369_reg            ;
wire [32-1:0] jump_type370_reg            ;
wire [32-1:0] jump_type371_reg            ;
wire [32-1:0] jump_type372_reg            ;
wire [32-1:0] jump_type373_reg            ;
wire [32-1:0] jump_type374_reg            ;
wire [32-1:0] jump_type375_reg            ;
wire [32-1:0] jump_type376_reg            ;
wire [32-1:0] jump_type377_reg            ;
wire [32-1:0] jump_type378_reg            ;
wire [32-1:0] jump_type379_reg            ;
wire [32-1:0] jump_type380_reg            ;
wire [32-1:0] jump_type381_reg            ;
wire [32-1:0] jump_type382_reg            ;
wire [32-1:0] jump_type383_reg            ;
wire [32-1:0] jump_type384_reg            ;
wire [32-1:0] jump_type385_reg            ;
wire [32-1:0] jump_type386_reg            ;
wire [32-1:0] jump_type387_reg            ;
wire [32-1:0] jump_type388_reg            ;
wire [32-1:0] jump_type389_reg            ;
wire [32-1:0] jump_type390_reg            ;
wire [32-1:0] jump_type391_reg            ;
wire [32-1:0] jump_type392_reg            ;
wire [32-1:0] jump_type393_reg            ;
wire [32-1:0] jump_type394_reg            ;
wire [32-1:0] jump_type395_reg            ;
wire [32-1:0] jump_type396_reg            ;
wire [32-1:0] jump_type397_reg            ;
wire [32-1:0] jump_type398_reg            ;
wire [32-1:0] jump_type399_reg            ;
wire [32-1:0] jump_type400_reg            ;
wire [32-1:0] jump_type401_reg            ;
wire [32-1:0] jump_type402_reg            ;
wire [32-1:0] jump_type403_reg            ;
wire [32-1:0] jump_type404_reg            ;
wire [32-1:0] jump_type405_reg            ;
wire [32-1:0] jump_type406_reg            ;
wire [32-1:0] jump_type407_reg            ;
wire [32-1:0] jump_type408_reg            ;
wire [32-1:0] jump_type409_reg            ;
wire [32-1:0] jump_type410_reg            ;
wire [32-1:0] jump_type411_reg            ;
wire [32-1:0] jump_type412_reg            ;
wire [32-1:0] jump_type413_reg            ;
wire [32-1:0] jump_type414_reg            ;
wire [32-1:0] jump_type415_reg            ;
wire [32-1:0] jump_type416_reg            ;
wire [32-1:0] jump_type417_reg            ;
wire [32-1:0] jump_type418_reg            ;
wire [32-1:0] jump_type419_reg            ;
wire [32-1:0] jump_type420_reg            ;
wire [32-1:0] jump_type421_reg            ;
wire [32-1:0] jump_type422_reg            ;
wire [32-1:0] jump_type423_reg            ;
wire [32-1:0] jump_type424_reg            ;
wire [32-1:0] jump_type425_reg            ;
wire [32-1:0] jump_type426_reg            ;
wire [32-1:0] jump_type427_reg            ;
wire [32-1:0] jump_type428_reg            ;
wire [32-1:0] jump_type429_reg            ;
wire [32-1:0] jump_type430_reg            ;
wire [32-1:0] jump_type431_reg            ;
wire [32-1:0] jump_type432_reg            ;
wire [32-1:0] jump_type433_reg            ;
wire [32-1:0] jump_type434_reg            ;
wire [32-1:0] jump_type435_reg            ;
wire [32-1:0] jump_type436_reg            ;
wire [32-1:0] jump_type437_reg            ;
wire [32-1:0] jump_type438_reg            ;
wire [32-1:0] jump_type439_reg            ;
wire [32-1:0] jump_type440_reg            ;
wire [32-1:0] jump_type441_reg            ;
wire [32-1:0] jump_type442_reg            ;
wire [32-1:0] jump_type443_reg            ;
wire [32-1:0] jump_type444_reg            ;
wire [32-1:0] jump_type445_reg            ;
wire [32-1:0] jump_type446_reg            ;
wire [32-1:0] jump_type447_reg            ;
wire [32-1:0] jump_type448_reg            ;
wire [32-1:0] jump_type449_reg            ;
wire [32-1:0] jump_type450_reg            ;
wire [32-1:0] jump_type451_reg            ;
wire [32-1:0] jump_type452_reg            ;
wire [32-1:0] jump_type453_reg            ;
wire [32-1:0] jump_type454_reg            ;
wire [32-1:0] jump_type455_reg            ;
wire [32-1:0] jump_type456_reg            ;
wire [32-1:0] jump_type457_reg            ;
wire [32-1:0] jump_type458_reg            ;
wire [32-1:0] jump_type459_reg            ;
wire [32-1:0] jump_type460_reg            ;
wire [32-1:0] jump_type461_reg            ;
wire [32-1:0] jump_type462_reg            ;
wire [32-1:0] jump_type463_reg            ;
wire [32-1:0] jump_type464_reg            ;
wire [32-1:0] jump_type465_reg            ;
wire [32-1:0] jump_type466_reg            ;
wire [32-1:0] jump_type467_reg            ;
wire [32-1:0] jump_type468_reg            ;
wire [32-1:0] jump_type469_reg            ;
wire [32-1:0] jump_type470_reg            ;
wire [32-1:0] jump_type471_reg            ;
wire [32-1:0] jump_type472_reg            ;
wire [32-1:0] jump_type473_reg            ;
wire [32-1:0] jump_type474_reg            ;
wire [32-1:0] jump_type475_reg            ;
wire [32-1:0] jump_type476_reg            ;
wire [32-1:0] jump_type477_reg            ;
wire [32-1:0] jump_type478_reg            ;
wire [32-1:0] jump_type479_reg            ;
wire [32-1:0] jump_type480_reg            ;
wire [32-1:0] jump_type481_reg            ;
wire [32-1:0] jump_type482_reg            ;
wire [32-1:0] jump_type483_reg            ;
wire [32-1:0] jump_type484_reg            ;
wire [32-1:0] jump_type485_reg            ;
wire [32-1:0] jump_type486_reg            ;
wire [32-1:0] jump_type487_reg            ;
wire [32-1:0] jump_type488_reg            ;
wire [32-1:0] jump_type489_reg            ;
wire [32-1:0] jump_type490_reg            ;
wire [32-1:0] jump_type491_reg            ;
wire [32-1:0] jump_type492_reg            ;
wire [32-1:0] jump_type493_reg            ;
wire [32-1:0] jump_type494_reg            ;
wire [32-1:0] jump_type495_reg            ;
wire [32-1:0] jump_type496_reg            ;
wire [32-1:0] jump_type497_reg            ;
wire [32-1:0] jump_type498_reg            ;
wire [32-1:0] jump_type499_reg            ;
wire [32-1:0] jump_type500_reg            ;
wire [32-1:0] jump_type501_reg            ;
wire [32-1:0] jump_type502_reg            ;
wire [32-1:0] jump_type503_reg            ;
wire [32-1:0] jump_type504_reg            ;
wire [32-1:0] jump_type505_reg            ;
wire [32-1:0] jump_type506_reg            ;
wire [32-1:0] jump_type507_reg            ;
wire [32-1:0] jump_type508_reg            ;
wire [32-1:0] jump_type509_reg            ;
wire [32-1:0] jump_type510_reg            ;
wire [32-1:0] jump_type511_reg            ;

//----------------------------control logic---------------------------------------------
wire common_para_wr               = ( waddr == COMMON_PARA_REG ) && wen;
wire jump_type0_wr                = ( waddr == JUMP_TYPE0_REG ) && wen;
wire jump_type1_wr                = ( waddr == JUMP_TYPE1_REG ) && wen;
wire jump_type2_wr                = ( waddr == JUMP_TYPE2_REG ) && wen;
wire jump_type3_wr                = ( waddr == JUMP_TYPE3_REG ) && wen;
wire jump_type4_wr                = ( waddr == JUMP_TYPE4_REG ) && wen;
wire jump_type5_wr                = ( waddr == JUMP_TYPE5_REG ) && wen;
wire jump_type6_wr                = ( waddr == JUMP_TYPE6_REG ) && wen;
wire jump_type7_wr                = ( waddr == JUMP_TYPE7_REG ) && wen;
wire jump_type8_wr                = ( waddr == JUMP_TYPE8_REG ) && wen;
wire jump_type9_wr                = ( waddr == JUMP_TYPE9_REG ) && wen;
wire jump_type10_wr               = ( waddr == JUMP_TYPE10_REG ) && wen;
wire jump_type11_wr               = ( waddr == JUMP_TYPE11_REG ) && wen;
wire jump_type12_wr               = ( waddr == JUMP_TYPE12_REG ) && wen;
wire jump_type13_wr               = ( waddr == JUMP_TYPE13_REG ) && wen;
wire jump_type14_wr               = ( waddr == JUMP_TYPE14_REG ) && wen;
wire jump_type15_wr               = ( waddr == JUMP_TYPE15_REG ) && wen;
wire jump_type16_wr               = ( waddr == JUMP_TYPE16_REG ) && wen;
wire jump_type17_wr               = ( waddr == JUMP_TYPE17_REG ) && wen;
wire jump_type18_wr               = ( waddr == JUMP_TYPE18_REG ) && wen;
wire jump_type19_wr               = ( waddr == JUMP_TYPE19_REG ) && wen;
wire jump_type20_wr               = ( waddr == JUMP_TYPE20_REG ) && wen;
wire jump_type21_wr               = ( waddr == JUMP_TYPE21_REG ) && wen;
wire jump_type22_wr               = ( waddr == JUMP_TYPE22_REG ) && wen;
wire jump_type23_wr               = ( waddr == JUMP_TYPE23_REG ) && wen;
wire jump_type24_wr               = ( waddr == JUMP_TYPE24_REG ) && wen;
wire jump_type25_wr               = ( waddr == JUMP_TYPE25_REG ) && wen;
wire jump_type26_wr               = ( waddr == JUMP_TYPE26_REG ) && wen;
wire jump_type27_wr               = ( waddr == JUMP_TYPE27_REG ) && wen;
wire jump_type28_wr               = ( waddr == JUMP_TYPE28_REG ) && wen;
wire jump_type29_wr               = ( waddr == JUMP_TYPE29_REG ) && wen;
wire jump_type30_wr               = ( waddr == JUMP_TYPE30_REG ) && wen;
wire jump_type31_wr               = ( waddr == JUMP_TYPE31_REG ) && wen;
wire jump_type32_wr               = ( waddr == JUMP_TYPE32_REG ) && wen;
wire jump_type33_wr               = ( waddr == JUMP_TYPE33_REG ) && wen;
wire jump_type34_wr               = ( waddr == JUMP_TYPE34_REG ) && wen;
wire jump_type35_wr               = ( waddr == JUMP_TYPE35_REG ) && wen;
wire jump_type36_wr               = ( waddr == JUMP_TYPE36_REG ) && wen;
wire jump_type37_wr               = ( waddr == JUMP_TYPE37_REG ) && wen;
wire jump_type38_wr               = ( waddr == JUMP_TYPE38_REG ) && wen;
wire jump_type39_wr               = ( waddr == JUMP_TYPE39_REG ) && wen;
wire jump_type40_wr               = ( waddr == JUMP_TYPE40_REG ) && wen;
wire jump_type41_wr               = ( waddr == JUMP_TYPE41_REG ) && wen;
wire jump_type42_wr               = ( waddr == JUMP_TYPE42_REG ) && wen;
wire jump_type43_wr               = ( waddr == JUMP_TYPE43_REG ) && wen;
wire jump_type44_wr               = ( waddr == JUMP_TYPE44_REG ) && wen;
wire jump_type45_wr               = ( waddr == JUMP_TYPE45_REG ) && wen;
wire jump_type46_wr               = ( waddr == JUMP_TYPE46_REG ) && wen;
wire jump_type47_wr               = ( waddr == JUMP_TYPE47_REG ) && wen;
wire jump_type48_wr               = ( waddr == JUMP_TYPE48_REG ) && wen;
wire jump_type49_wr               = ( waddr == JUMP_TYPE49_REG ) && wen;
wire jump_type50_wr               = ( waddr == JUMP_TYPE50_REG ) && wen;
wire jump_type51_wr               = ( waddr == JUMP_TYPE51_REG ) && wen;
wire jump_type52_wr               = ( waddr == JUMP_TYPE52_REG ) && wen;
wire jump_type53_wr               = ( waddr == JUMP_TYPE53_REG ) && wen;
wire jump_type54_wr               = ( waddr == JUMP_TYPE54_REG ) && wen;
wire jump_type55_wr               = ( waddr == JUMP_TYPE55_REG ) && wen;
wire jump_type56_wr               = ( waddr == JUMP_TYPE56_REG ) && wen;
wire jump_type57_wr               = ( waddr == JUMP_TYPE57_REG ) && wen;
wire jump_type58_wr               = ( waddr == JUMP_TYPE58_REG ) && wen;
wire jump_type59_wr               = ( waddr == JUMP_TYPE59_REG ) && wen;
wire jump_type60_wr               = ( waddr == JUMP_TYPE60_REG ) && wen;
wire jump_type61_wr               = ( waddr == JUMP_TYPE61_REG ) && wen;
wire jump_type62_wr               = ( waddr == JUMP_TYPE62_REG ) && wen;
wire jump_type63_wr               = ( waddr == JUMP_TYPE63_REG ) && wen;
wire jump_type64_wr               = ( waddr == JUMP_TYPE64_REG ) && wen;
wire jump_type65_wr               = ( waddr == JUMP_TYPE65_REG ) && wen;
wire jump_type66_wr               = ( waddr == JUMP_TYPE66_REG ) && wen;
wire jump_type67_wr               = ( waddr == JUMP_TYPE67_REG ) && wen;
wire jump_type68_wr               = ( waddr == JUMP_TYPE68_REG ) && wen;
wire jump_type69_wr               = ( waddr == JUMP_TYPE69_REG ) && wen;
wire jump_type70_wr               = ( waddr == JUMP_TYPE70_REG ) && wen;
wire jump_type71_wr               = ( waddr == JUMP_TYPE71_REG ) && wen;
wire jump_type72_wr               = ( waddr == JUMP_TYPE72_REG ) && wen;
wire jump_type73_wr               = ( waddr == JUMP_TYPE73_REG ) && wen;
wire jump_type74_wr               = ( waddr == JUMP_TYPE74_REG ) && wen;
wire jump_type75_wr               = ( waddr == JUMP_TYPE75_REG ) && wen;
wire jump_type76_wr               = ( waddr == JUMP_TYPE76_REG ) && wen;
wire jump_type77_wr               = ( waddr == JUMP_TYPE77_REG ) && wen;
wire jump_type78_wr               = ( waddr == JUMP_TYPE78_REG ) && wen;
wire jump_type79_wr               = ( waddr == JUMP_TYPE79_REG ) && wen;
wire jump_type80_wr               = ( waddr == JUMP_TYPE80_REG ) && wen;
wire jump_type81_wr               = ( waddr == JUMP_TYPE81_REG ) && wen;
wire jump_type82_wr               = ( waddr == JUMP_TYPE82_REG ) && wen;
wire jump_type83_wr               = ( waddr == JUMP_TYPE83_REG ) && wen;
wire jump_type84_wr               = ( waddr == JUMP_TYPE84_REG ) && wen;
wire jump_type85_wr               = ( waddr == JUMP_TYPE85_REG ) && wen;
wire jump_type86_wr               = ( waddr == JUMP_TYPE86_REG ) && wen;
wire jump_type87_wr               = ( waddr == JUMP_TYPE87_REG ) && wen;
wire jump_type88_wr               = ( waddr == JUMP_TYPE88_REG ) && wen;
wire jump_type89_wr               = ( waddr == JUMP_TYPE89_REG ) && wen;
wire jump_type90_wr               = ( waddr == JUMP_TYPE90_REG ) && wen;
wire jump_type91_wr               = ( waddr == JUMP_TYPE91_REG ) && wen;
wire jump_type92_wr               = ( waddr == JUMP_TYPE92_REG ) && wen;
wire jump_type93_wr               = ( waddr == JUMP_TYPE93_REG ) && wen;
wire jump_type94_wr               = ( waddr == JUMP_TYPE94_REG ) && wen;
wire jump_type95_wr               = ( waddr == JUMP_TYPE95_REG ) && wen;
wire jump_type96_wr               = ( waddr == JUMP_TYPE96_REG ) && wen;
wire jump_type97_wr               = ( waddr == JUMP_TYPE97_REG ) && wen;
wire jump_type98_wr               = ( waddr == JUMP_TYPE98_REG ) && wen;
wire jump_type99_wr               = ( waddr == JUMP_TYPE99_REG ) && wen;
wire jump_type100_wr              = ( waddr == JUMP_TYPE100_REG ) && wen;
wire jump_type101_wr              = ( waddr == JUMP_TYPE101_REG ) && wen;
wire jump_type102_wr              = ( waddr == JUMP_TYPE102_REG ) && wen;
wire jump_type103_wr              = ( waddr == JUMP_TYPE103_REG ) && wen;
wire jump_type104_wr              = ( waddr == JUMP_TYPE104_REG ) && wen;
wire jump_type105_wr              = ( waddr == JUMP_TYPE105_REG ) && wen;
wire jump_type106_wr              = ( waddr == JUMP_TYPE106_REG ) && wen;
wire jump_type107_wr              = ( waddr == JUMP_TYPE107_REG ) && wen;
wire jump_type108_wr              = ( waddr == JUMP_TYPE108_REG ) && wen;
wire jump_type109_wr              = ( waddr == JUMP_TYPE109_REG ) && wen;
wire jump_type110_wr              = ( waddr == JUMP_TYPE110_REG ) && wen;
wire jump_type111_wr              = ( waddr == JUMP_TYPE111_REG ) && wen;
wire jump_type112_wr              = ( waddr == JUMP_TYPE112_REG ) && wen;
wire jump_type113_wr              = ( waddr == JUMP_TYPE113_REG ) && wen;
wire jump_type114_wr              = ( waddr == JUMP_TYPE114_REG ) && wen;
wire jump_type115_wr              = ( waddr == JUMP_TYPE115_REG ) && wen;
wire jump_type116_wr              = ( waddr == JUMP_TYPE116_REG ) && wen;
wire jump_type117_wr              = ( waddr == JUMP_TYPE117_REG ) && wen;
wire jump_type118_wr              = ( waddr == JUMP_TYPE118_REG ) && wen;
wire jump_type119_wr              = ( waddr == JUMP_TYPE119_REG ) && wen;
wire jump_type120_wr              = ( waddr == JUMP_TYPE120_REG ) && wen;
wire jump_type121_wr              = ( waddr == JUMP_TYPE121_REG ) && wen;
wire jump_type122_wr              = ( waddr == JUMP_TYPE122_REG ) && wen;
wire jump_type123_wr              = ( waddr == JUMP_TYPE123_REG ) && wen;
wire jump_type124_wr              = ( waddr == JUMP_TYPE124_REG ) && wen;
wire jump_type125_wr              = ( waddr == JUMP_TYPE125_REG ) && wen;
wire jump_type126_wr              = ( waddr == JUMP_TYPE126_REG ) && wen;
wire jump_type127_wr              = ( waddr == JUMP_TYPE127_REG ) && wen;
wire jump_type128_wr              = ( waddr == JUMP_TYPE128_REG ) && wen;
wire jump_type129_wr              = ( waddr == JUMP_TYPE129_REG ) && wen;
wire jump_type130_wr              = ( waddr == JUMP_TYPE130_REG ) && wen;
wire jump_type131_wr              = ( waddr == JUMP_TYPE131_REG ) && wen;
wire jump_type132_wr              = ( waddr == JUMP_TYPE132_REG ) && wen;
wire jump_type133_wr              = ( waddr == JUMP_TYPE133_REG ) && wen;
wire jump_type134_wr              = ( waddr == JUMP_TYPE134_REG ) && wen;
wire jump_type135_wr              = ( waddr == JUMP_TYPE135_REG ) && wen;
wire jump_type136_wr              = ( waddr == JUMP_TYPE136_REG ) && wen;
wire jump_type137_wr              = ( waddr == JUMP_TYPE137_REG ) && wen;
wire jump_type138_wr              = ( waddr == JUMP_TYPE138_REG ) && wen;
wire jump_type139_wr              = ( waddr == JUMP_TYPE139_REG ) && wen;
wire jump_type140_wr              = ( waddr == JUMP_TYPE140_REG ) && wen;
wire jump_type141_wr              = ( waddr == JUMP_TYPE141_REG ) && wen;
wire jump_type142_wr              = ( waddr == JUMP_TYPE142_REG ) && wen;
wire jump_type143_wr              = ( waddr == JUMP_TYPE143_REG ) && wen;
wire jump_type144_wr              = ( waddr == JUMP_TYPE144_REG ) && wen;
wire jump_type145_wr              = ( waddr == JUMP_TYPE145_REG ) && wen;
wire jump_type146_wr              = ( waddr == JUMP_TYPE146_REG ) && wen;
wire jump_type147_wr              = ( waddr == JUMP_TYPE147_REG ) && wen;
wire jump_type148_wr              = ( waddr == JUMP_TYPE148_REG ) && wen;
wire jump_type149_wr              = ( waddr == JUMP_TYPE149_REG ) && wen;
wire jump_type150_wr              = ( waddr == JUMP_TYPE150_REG ) && wen;
wire jump_type151_wr              = ( waddr == JUMP_TYPE151_REG ) && wen;
wire jump_type152_wr              = ( waddr == JUMP_TYPE152_REG ) && wen;
wire jump_type153_wr              = ( waddr == JUMP_TYPE153_REG ) && wen;
wire jump_type154_wr              = ( waddr == JUMP_TYPE154_REG ) && wen;
wire jump_type155_wr              = ( waddr == JUMP_TYPE155_REG ) && wen;
wire jump_type156_wr              = ( waddr == JUMP_TYPE156_REG ) && wen;
wire jump_type157_wr              = ( waddr == JUMP_TYPE157_REG ) && wen;
wire jump_type158_wr              = ( waddr == JUMP_TYPE158_REG ) && wen;
wire jump_type159_wr              = ( waddr == JUMP_TYPE159_REG ) && wen;
wire jump_type160_wr              = ( waddr == JUMP_TYPE160_REG ) && wen;
wire jump_type161_wr              = ( waddr == JUMP_TYPE161_REG ) && wen;
wire jump_type162_wr              = ( waddr == JUMP_TYPE162_REG ) && wen;
wire jump_type163_wr              = ( waddr == JUMP_TYPE163_REG ) && wen;
wire jump_type164_wr              = ( waddr == JUMP_TYPE164_REG ) && wen;
wire jump_type165_wr              = ( waddr == JUMP_TYPE165_REG ) && wen;
wire jump_type166_wr              = ( waddr == JUMP_TYPE166_REG ) && wen;
wire jump_type167_wr              = ( waddr == JUMP_TYPE167_REG ) && wen;
wire jump_type168_wr              = ( waddr == JUMP_TYPE168_REG ) && wen;
wire jump_type169_wr              = ( waddr == JUMP_TYPE169_REG ) && wen;
wire jump_type170_wr              = ( waddr == JUMP_TYPE170_REG ) && wen;
wire jump_type171_wr              = ( waddr == JUMP_TYPE171_REG ) && wen;
wire jump_type172_wr              = ( waddr == JUMP_TYPE172_REG ) && wen;
wire jump_type173_wr              = ( waddr == JUMP_TYPE173_REG ) && wen;
wire jump_type174_wr              = ( waddr == JUMP_TYPE174_REG ) && wen;
wire jump_type175_wr              = ( waddr == JUMP_TYPE175_REG ) && wen;
wire jump_type176_wr              = ( waddr == JUMP_TYPE176_REG ) && wen;
wire jump_type177_wr              = ( waddr == JUMP_TYPE177_REG ) && wen;
wire jump_type178_wr              = ( waddr == JUMP_TYPE178_REG ) && wen;
wire jump_type179_wr              = ( waddr == JUMP_TYPE179_REG ) && wen;
wire jump_type180_wr              = ( waddr == JUMP_TYPE180_REG ) && wen;
wire jump_type181_wr              = ( waddr == JUMP_TYPE181_REG ) && wen;
wire jump_type182_wr              = ( waddr == JUMP_TYPE182_REG ) && wen;
wire jump_type183_wr              = ( waddr == JUMP_TYPE183_REG ) && wen;
wire jump_type184_wr              = ( waddr == JUMP_TYPE184_REG ) && wen;
wire jump_type185_wr              = ( waddr == JUMP_TYPE185_REG ) && wen;
wire jump_type186_wr              = ( waddr == JUMP_TYPE186_REG ) && wen;
wire jump_type187_wr              = ( waddr == JUMP_TYPE187_REG ) && wen;
wire jump_type188_wr              = ( waddr == JUMP_TYPE188_REG ) && wen;
wire jump_type189_wr              = ( waddr == JUMP_TYPE189_REG ) && wen;
wire jump_type190_wr              = ( waddr == JUMP_TYPE190_REG ) && wen;
wire jump_type191_wr              = ( waddr == JUMP_TYPE191_REG ) && wen;
wire jump_type192_wr              = ( waddr == JUMP_TYPE192_REG ) && wen;
wire jump_type193_wr              = ( waddr == JUMP_TYPE193_REG ) && wen;
wire jump_type194_wr              = ( waddr == JUMP_TYPE194_REG ) && wen;
wire jump_type195_wr              = ( waddr == JUMP_TYPE195_REG ) && wen;
wire jump_type196_wr              = ( waddr == JUMP_TYPE196_REG ) && wen;
wire jump_type197_wr              = ( waddr == JUMP_TYPE197_REG ) && wen;
wire jump_type198_wr              = ( waddr == JUMP_TYPE198_REG ) && wen;
wire jump_type199_wr              = ( waddr == JUMP_TYPE199_REG ) && wen;
wire jump_type200_wr              = ( waddr == JUMP_TYPE200_REG ) && wen;
wire jump_type201_wr              = ( waddr == JUMP_TYPE201_REG ) && wen;
wire jump_type202_wr              = ( waddr == JUMP_TYPE202_REG ) && wen;
wire jump_type203_wr              = ( waddr == JUMP_TYPE203_REG ) && wen;
wire jump_type204_wr              = ( waddr == JUMP_TYPE204_REG ) && wen;
wire jump_type205_wr              = ( waddr == JUMP_TYPE205_REG ) && wen;
wire jump_type206_wr              = ( waddr == JUMP_TYPE206_REG ) && wen;
wire jump_type207_wr              = ( waddr == JUMP_TYPE207_REG ) && wen;
wire jump_type208_wr              = ( waddr == JUMP_TYPE208_REG ) && wen;
wire jump_type209_wr              = ( waddr == JUMP_TYPE209_REG ) && wen;
wire jump_type210_wr              = ( waddr == JUMP_TYPE210_REG ) && wen;
wire jump_type211_wr              = ( waddr == JUMP_TYPE211_REG ) && wen;
wire jump_type212_wr              = ( waddr == JUMP_TYPE212_REG ) && wen;
wire jump_type213_wr              = ( waddr == JUMP_TYPE213_REG ) && wen;
wire jump_type214_wr              = ( waddr == JUMP_TYPE214_REG ) && wen;
wire jump_type215_wr              = ( waddr == JUMP_TYPE215_REG ) && wen;
wire jump_type216_wr              = ( waddr == JUMP_TYPE216_REG ) && wen;
wire jump_type217_wr              = ( waddr == JUMP_TYPE217_REG ) && wen;
wire jump_type218_wr              = ( waddr == JUMP_TYPE218_REG ) && wen;
wire jump_type219_wr              = ( waddr == JUMP_TYPE219_REG ) && wen;
wire jump_type220_wr              = ( waddr == JUMP_TYPE220_REG ) && wen;
wire jump_type221_wr              = ( waddr == JUMP_TYPE221_REG ) && wen;
wire jump_type222_wr              = ( waddr == JUMP_TYPE222_REG ) && wen;
wire jump_type223_wr              = ( waddr == JUMP_TYPE223_REG ) && wen;
wire jump_type224_wr              = ( waddr == JUMP_TYPE224_REG ) && wen;
wire jump_type225_wr              = ( waddr == JUMP_TYPE225_REG ) && wen;
wire jump_type226_wr              = ( waddr == JUMP_TYPE226_REG ) && wen;
wire jump_type227_wr              = ( waddr == JUMP_TYPE227_REG ) && wen;
wire jump_type228_wr              = ( waddr == JUMP_TYPE228_REG ) && wen;
wire jump_type229_wr              = ( waddr == JUMP_TYPE229_REG ) && wen;
wire jump_type230_wr              = ( waddr == JUMP_TYPE230_REG ) && wen;
wire jump_type231_wr              = ( waddr == JUMP_TYPE231_REG ) && wen;
wire jump_type232_wr              = ( waddr == JUMP_TYPE232_REG ) && wen;
wire jump_type233_wr              = ( waddr == JUMP_TYPE233_REG ) && wen;
wire jump_type234_wr              = ( waddr == JUMP_TYPE234_REG ) && wen;
wire jump_type235_wr              = ( waddr == JUMP_TYPE235_REG ) && wen;
wire jump_type236_wr              = ( waddr == JUMP_TYPE236_REG ) && wen;
wire jump_type237_wr              = ( waddr == JUMP_TYPE237_REG ) && wen;
wire jump_type238_wr              = ( waddr == JUMP_TYPE238_REG ) && wen;
wire jump_type239_wr              = ( waddr == JUMP_TYPE239_REG ) && wen;
wire jump_type240_wr              = ( waddr == JUMP_TYPE240_REG ) && wen;
wire jump_type241_wr              = ( waddr == JUMP_TYPE241_REG ) && wen;
wire jump_type242_wr              = ( waddr == JUMP_TYPE242_REG ) && wen;
wire jump_type243_wr              = ( waddr == JUMP_TYPE243_REG ) && wen;
wire jump_type244_wr              = ( waddr == JUMP_TYPE244_REG ) && wen;
wire jump_type245_wr              = ( waddr == JUMP_TYPE245_REG ) && wen;
wire jump_type246_wr              = ( waddr == JUMP_TYPE246_REG ) && wen;
wire jump_type247_wr              = ( waddr == JUMP_TYPE247_REG ) && wen;
wire jump_type248_wr              = ( waddr == JUMP_TYPE248_REG ) && wen;
wire jump_type249_wr              = ( waddr == JUMP_TYPE249_REG ) && wen;
wire jump_type250_wr              = ( waddr == JUMP_TYPE250_REG ) && wen;
wire jump_type251_wr              = ( waddr == JUMP_TYPE251_REG ) && wen;
wire jump_type252_wr              = ( waddr == JUMP_TYPE252_REG ) && wen;
wire jump_type253_wr              = ( waddr == JUMP_TYPE253_REG ) && wen;
wire jump_type254_wr              = ( waddr == JUMP_TYPE254_REG ) && wen;
wire jump_type255_wr              = ( waddr == JUMP_TYPE255_REG ) && wen;
wire jump_type256_wr              = ( waddr == JUMP_TYPE256_REG ) && wen;
wire jump_type257_wr              = ( waddr == JUMP_TYPE257_REG ) && wen;
wire jump_type258_wr              = ( waddr == JUMP_TYPE258_REG ) && wen;
wire jump_type259_wr              = ( waddr == JUMP_TYPE259_REG ) && wen;
wire jump_type260_wr              = ( waddr == JUMP_TYPE260_REG ) && wen;
wire jump_type261_wr              = ( waddr == JUMP_TYPE261_REG ) && wen;
wire jump_type262_wr              = ( waddr == JUMP_TYPE262_REG ) && wen;
wire jump_type263_wr              = ( waddr == JUMP_TYPE263_REG ) && wen;
wire jump_type264_wr              = ( waddr == JUMP_TYPE264_REG ) && wen;
wire jump_type265_wr              = ( waddr == JUMP_TYPE265_REG ) && wen;
wire jump_type266_wr              = ( waddr == JUMP_TYPE266_REG ) && wen;
wire jump_type267_wr              = ( waddr == JUMP_TYPE267_REG ) && wen;
wire jump_type268_wr              = ( waddr == JUMP_TYPE268_REG ) && wen;
wire jump_type269_wr              = ( waddr == JUMP_TYPE269_REG ) && wen;
wire jump_type270_wr              = ( waddr == JUMP_TYPE270_REG ) && wen;
wire jump_type271_wr              = ( waddr == JUMP_TYPE271_REG ) && wen;
wire jump_type272_wr              = ( waddr == JUMP_TYPE272_REG ) && wen;
wire jump_type273_wr              = ( waddr == JUMP_TYPE273_REG ) && wen;
wire jump_type274_wr              = ( waddr == JUMP_TYPE274_REG ) && wen;
wire jump_type275_wr              = ( waddr == JUMP_TYPE275_REG ) && wen;
wire jump_type276_wr              = ( waddr == JUMP_TYPE276_REG ) && wen;
wire jump_type277_wr              = ( waddr == JUMP_TYPE277_REG ) && wen;
wire jump_type278_wr              = ( waddr == JUMP_TYPE278_REG ) && wen;
wire jump_type279_wr              = ( waddr == JUMP_TYPE279_REG ) && wen;
wire jump_type280_wr              = ( waddr == JUMP_TYPE280_REG ) && wen;
wire jump_type281_wr              = ( waddr == JUMP_TYPE281_REG ) && wen;
wire jump_type282_wr              = ( waddr == JUMP_TYPE282_REG ) && wen;
wire jump_type283_wr              = ( waddr == JUMP_TYPE283_REG ) && wen;
wire jump_type284_wr              = ( waddr == JUMP_TYPE284_REG ) && wen;
wire jump_type285_wr              = ( waddr == JUMP_TYPE285_REG ) && wen;
wire jump_type286_wr              = ( waddr == JUMP_TYPE286_REG ) && wen;
wire jump_type287_wr              = ( waddr == JUMP_TYPE287_REG ) && wen;
wire jump_type288_wr              = ( waddr == JUMP_TYPE288_REG ) && wen;
wire jump_type289_wr              = ( waddr == JUMP_TYPE289_REG ) && wen;
wire jump_type290_wr              = ( waddr == JUMP_TYPE290_REG ) && wen;
wire jump_type291_wr              = ( waddr == JUMP_TYPE291_REG ) && wen;
wire jump_type292_wr              = ( waddr == JUMP_TYPE292_REG ) && wen;
wire jump_type293_wr              = ( waddr == JUMP_TYPE293_REG ) && wen;
wire jump_type294_wr              = ( waddr == JUMP_TYPE294_REG ) && wen;
wire jump_type295_wr              = ( waddr == JUMP_TYPE295_REG ) && wen;
wire jump_type296_wr              = ( waddr == JUMP_TYPE296_REG ) && wen;
wire jump_type297_wr              = ( waddr == JUMP_TYPE297_REG ) && wen;
wire jump_type298_wr              = ( waddr == JUMP_TYPE298_REG ) && wen;
wire jump_type299_wr              = ( waddr == JUMP_TYPE299_REG ) && wen;
wire jump_type300_wr              = ( waddr == JUMP_TYPE300_REG ) && wen;
wire jump_type301_wr              = ( waddr == JUMP_TYPE301_REG ) && wen;
wire jump_type302_wr              = ( waddr == JUMP_TYPE302_REG ) && wen;
wire jump_type303_wr              = ( waddr == JUMP_TYPE303_REG ) && wen;
wire jump_type304_wr              = ( waddr == JUMP_TYPE304_REG ) && wen;
wire jump_type305_wr              = ( waddr == JUMP_TYPE305_REG ) && wen;
wire jump_type306_wr              = ( waddr == JUMP_TYPE306_REG ) && wen;
wire jump_type307_wr              = ( waddr == JUMP_TYPE307_REG ) && wen;
wire jump_type308_wr              = ( waddr == JUMP_TYPE308_REG ) && wen;
wire jump_type309_wr              = ( waddr == JUMP_TYPE309_REG ) && wen;
wire jump_type310_wr              = ( waddr == JUMP_TYPE310_REG ) && wen;
wire jump_type311_wr              = ( waddr == JUMP_TYPE311_REG ) && wen;
wire jump_type312_wr              = ( waddr == JUMP_TYPE312_REG ) && wen;
wire jump_type313_wr              = ( waddr == JUMP_TYPE313_REG ) && wen;
wire jump_type314_wr              = ( waddr == JUMP_TYPE314_REG ) && wen;
wire jump_type315_wr              = ( waddr == JUMP_TYPE315_REG ) && wen;
wire jump_type316_wr              = ( waddr == JUMP_TYPE316_REG ) && wen;
wire jump_type317_wr              = ( waddr == JUMP_TYPE317_REG ) && wen;
wire jump_type318_wr              = ( waddr == JUMP_TYPE318_REG ) && wen;
wire jump_type319_wr              = ( waddr == JUMP_TYPE319_REG ) && wen;
wire jump_type320_wr              = ( waddr == JUMP_TYPE320_REG ) && wen;
wire jump_type321_wr              = ( waddr == JUMP_TYPE321_REG ) && wen;
wire jump_type322_wr              = ( waddr == JUMP_TYPE322_REG ) && wen;
wire jump_type323_wr              = ( waddr == JUMP_TYPE323_REG ) && wen;
wire jump_type324_wr              = ( waddr == JUMP_TYPE324_REG ) && wen;
wire jump_type325_wr              = ( waddr == JUMP_TYPE325_REG ) && wen;
wire jump_type326_wr              = ( waddr == JUMP_TYPE326_REG ) && wen;
wire jump_type327_wr              = ( waddr == JUMP_TYPE327_REG ) && wen;
wire jump_type328_wr              = ( waddr == JUMP_TYPE328_REG ) && wen;
wire jump_type329_wr              = ( waddr == JUMP_TYPE329_REG ) && wen;
wire jump_type330_wr              = ( waddr == JUMP_TYPE330_REG ) && wen;
wire jump_type331_wr              = ( waddr == JUMP_TYPE331_REG ) && wen;
wire jump_type332_wr              = ( waddr == JUMP_TYPE332_REG ) && wen;
wire jump_type333_wr              = ( waddr == JUMP_TYPE333_REG ) && wen;
wire jump_type334_wr              = ( waddr == JUMP_TYPE334_REG ) && wen;
wire jump_type335_wr              = ( waddr == JUMP_TYPE335_REG ) && wen;
wire jump_type336_wr              = ( waddr == JUMP_TYPE336_REG ) && wen;
wire jump_type337_wr              = ( waddr == JUMP_TYPE337_REG ) && wen;
wire jump_type338_wr              = ( waddr == JUMP_TYPE338_REG ) && wen;
wire jump_type339_wr              = ( waddr == JUMP_TYPE339_REG ) && wen;
wire jump_type340_wr              = ( waddr == JUMP_TYPE340_REG ) && wen;
wire jump_type341_wr              = ( waddr == JUMP_TYPE341_REG ) && wen;
wire jump_type342_wr              = ( waddr == JUMP_TYPE342_REG ) && wen;
wire jump_type343_wr              = ( waddr == JUMP_TYPE343_REG ) && wen;
wire jump_type344_wr              = ( waddr == JUMP_TYPE344_REG ) && wen;
wire jump_type345_wr              = ( waddr == JUMP_TYPE345_REG ) && wen;
wire jump_type346_wr              = ( waddr == JUMP_TYPE346_REG ) && wen;
wire jump_type347_wr              = ( waddr == JUMP_TYPE347_REG ) && wen;
wire jump_type348_wr              = ( waddr == JUMP_TYPE348_REG ) && wen;
wire jump_type349_wr              = ( waddr == JUMP_TYPE349_REG ) && wen;
wire jump_type350_wr              = ( waddr == JUMP_TYPE350_REG ) && wen;
wire jump_type351_wr              = ( waddr == JUMP_TYPE351_REG ) && wen;
wire jump_type352_wr              = ( waddr == JUMP_TYPE352_REG ) && wen;
wire jump_type353_wr              = ( waddr == JUMP_TYPE353_REG ) && wen;
wire jump_type354_wr              = ( waddr == JUMP_TYPE354_REG ) && wen;
wire jump_type355_wr              = ( waddr == JUMP_TYPE355_REG ) && wen;
wire jump_type356_wr              = ( waddr == JUMP_TYPE356_REG ) && wen;
wire jump_type357_wr              = ( waddr == JUMP_TYPE357_REG ) && wen;
wire jump_type358_wr              = ( waddr == JUMP_TYPE358_REG ) && wen;
wire jump_type359_wr              = ( waddr == JUMP_TYPE359_REG ) && wen;
wire jump_type360_wr              = ( waddr == JUMP_TYPE360_REG ) && wen;
wire jump_type361_wr              = ( waddr == JUMP_TYPE361_REG ) && wen;
wire jump_type362_wr              = ( waddr == JUMP_TYPE362_REG ) && wen;
wire jump_type363_wr              = ( waddr == JUMP_TYPE363_REG ) && wen;
wire jump_type364_wr              = ( waddr == JUMP_TYPE364_REG ) && wen;
wire jump_type365_wr              = ( waddr == JUMP_TYPE365_REG ) && wen;
wire jump_type366_wr              = ( waddr == JUMP_TYPE366_REG ) && wen;
wire jump_type367_wr              = ( waddr == JUMP_TYPE367_REG ) && wen;
wire jump_type368_wr              = ( waddr == JUMP_TYPE368_REG ) && wen;
wire jump_type369_wr              = ( waddr == JUMP_TYPE369_REG ) && wen;
wire jump_type370_wr              = ( waddr == JUMP_TYPE370_REG ) && wen;
wire jump_type371_wr              = ( waddr == JUMP_TYPE371_REG ) && wen;
wire jump_type372_wr              = ( waddr == JUMP_TYPE372_REG ) && wen;
wire jump_type373_wr              = ( waddr == JUMP_TYPE373_REG ) && wen;
wire jump_type374_wr              = ( waddr == JUMP_TYPE374_REG ) && wen;
wire jump_type375_wr              = ( waddr == JUMP_TYPE375_REG ) && wen;
wire jump_type376_wr              = ( waddr == JUMP_TYPE376_REG ) && wen;
wire jump_type377_wr              = ( waddr == JUMP_TYPE377_REG ) && wen;
wire jump_type378_wr              = ( waddr == JUMP_TYPE378_REG ) && wen;
wire jump_type379_wr              = ( waddr == JUMP_TYPE379_REG ) && wen;
wire jump_type380_wr              = ( waddr == JUMP_TYPE380_REG ) && wen;
wire jump_type381_wr              = ( waddr == JUMP_TYPE381_REG ) && wen;
wire jump_type382_wr              = ( waddr == JUMP_TYPE382_REG ) && wen;
wire jump_type383_wr              = ( waddr == JUMP_TYPE383_REG ) && wen;
wire jump_type384_wr              = ( waddr == JUMP_TYPE384_REG ) && wen;
wire jump_type385_wr              = ( waddr == JUMP_TYPE385_REG ) && wen;
wire jump_type386_wr              = ( waddr == JUMP_TYPE386_REG ) && wen;
wire jump_type387_wr              = ( waddr == JUMP_TYPE387_REG ) && wen;
wire jump_type388_wr              = ( waddr == JUMP_TYPE388_REG ) && wen;
wire jump_type389_wr              = ( waddr == JUMP_TYPE389_REG ) && wen;
wire jump_type390_wr              = ( waddr == JUMP_TYPE390_REG ) && wen;
wire jump_type391_wr              = ( waddr == JUMP_TYPE391_REG ) && wen;
wire jump_type392_wr              = ( waddr == JUMP_TYPE392_REG ) && wen;
wire jump_type393_wr              = ( waddr == JUMP_TYPE393_REG ) && wen;
wire jump_type394_wr              = ( waddr == JUMP_TYPE394_REG ) && wen;
wire jump_type395_wr              = ( waddr == JUMP_TYPE395_REG ) && wen;
wire jump_type396_wr              = ( waddr == JUMP_TYPE396_REG ) && wen;
wire jump_type397_wr              = ( waddr == JUMP_TYPE397_REG ) && wen;
wire jump_type398_wr              = ( waddr == JUMP_TYPE398_REG ) && wen;
wire jump_type399_wr              = ( waddr == JUMP_TYPE399_REG ) && wen;
wire jump_type400_wr              = ( waddr == JUMP_TYPE400_REG ) && wen;
wire jump_type401_wr              = ( waddr == JUMP_TYPE401_REG ) && wen;
wire jump_type402_wr              = ( waddr == JUMP_TYPE402_REG ) && wen;
wire jump_type403_wr              = ( waddr == JUMP_TYPE403_REG ) && wen;
wire jump_type404_wr              = ( waddr == JUMP_TYPE404_REG ) && wen;
wire jump_type405_wr              = ( waddr == JUMP_TYPE405_REG ) && wen;
wire jump_type406_wr              = ( waddr == JUMP_TYPE406_REG ) && wen;
wire jump_type407_wr              = ( waddr == JUMP_TYPE407_REG ) && wen;
wire jump_type408_wr              = ( waddr == JUMP_TYPE408_REG ) && wen;
wire jump_type409_wr              = ( waddr == JUMP_TYPE409_REG ) && wen;
wire jump_type410_wr              = ( waddr == JUMP_TYPE410_REG ) && wen;
wire jump_type411_wr              = ( waddr == JUMP_TYPE411_REG ) && wen;
wire jump_type412_wr              = ( waddr == JUMP_TYPE412_REG ) && wen;
wire jump_type413_wr              = ( waddr == JUMP_TYPE413_REG ) && wen;
wire jump_type414_wr              = ( waddr == JUMP_TYPE414_REG ) && wen;
wire jump_type415_wr              = ( waddr == JUMP_TYPE415_REG ) && wen;
wire jump_type416_wr              = ( waddr == JUMP_TYPE416_REG ) && wen;
wire jump_type417_wr              = ( waddr == JUMP_TYPE417_REG ) && wen;
wire jump_type418_wr              = ( waddr == JUMP_TYPE418_REG ) && wen;
wire jump_type419_wr              = ( waddr == JUMP_TYPE419_REG ) && wen;
wire jump_type420_wr              = ( waddr == JUMP_TYPE420_REG ) && wen;
wire jump_type421_wr              = ( waddr == JUMP_TYPE421_REG ) && wen;
wire jump_type422_wr              = ( waddr == JUMP_TYPE422_REG ) && wen;
wire jump_type423_wr              = ( waddr == JUMP_TYPE423_REG ) && wen;
wire jump_type424_wr              = ( waddr == JUMP_TYPE424_REG ) && wen;
wire jump_type425_wr              = ( waddr == JUMP_TYPE425_REG ) && wen;
wire jump_type426_wr              = ( waddr == JUMP_TYPE426_REG ) && wen;
wire jump_type427_wr              = ( waddr == JUMP_TYPE427_REG ) && wen;
wire jump_type428_wr              = ( waddr == JUMP_TYPE428_REG ) && wen;
wire jump_type429_wr              = ( waddr == JUMP_TYPE429_REG ) && wen;
wire jump_type430_wr              = ( waddr == JUMP_TYPE430_REG ) && wen;
wire jump_type431_wr              = ( waddr == JUMP_TYPE431_REG ) && wen;
wire jump_type432_wr              = ( waddr == JUMP_TYPE432_REG ) && wen;
wire jump_type433_wr              = ( waddr == JUMP_TYPE433_REG ) && wen;
wire jump_type434_wr              = ( waddr == JUMP_TYPE434_REG ) && wen;
wire jump_type435_wr              = ( waddr == JUMP_TYPE435_REG ) && wen;
wire jump_type436_wr              = ( waddr == JUMP_TYPE436_REG ) && wen;
wire jump_type437_wr              = ( waddr == JUMP_TYPE437_REG ) && wen;
wire jump_type438_wr              = ( waddr == JUMP_TYPE438_REG ) && wen;
wire jump_type439_wr              = ( waddr == JUMP_TYPE439_REG ) && wen;
wire jump_type440_wr              = ( waddr == JUMP_TYPE440_REG ) && wen;
wire jump_type441_wr              = ( waddr == JUMP_TYPE441_REG ) && wen;
wire jump_type442_wr              = ( waddr == JUMP_TYPE442_REG ) && wen;
wire jump_type443_wr              = ( waddr == JUMP_TYPE443_REG ) && wen;
wire jump_type444_wr              = ( waddr == JUMP_TYPE444_REG ) && wen;
wire jump_type445_wr              = ( waddr == JUMP_TYPE445_REG ) && wen;
wire jump_type446_wr              = ( waddr == JUMP_TYPE446_REG ) && wen;
wire jump_type447_wr              = ( waddr == JUMP_TYPE447_REG ) && wen;
wire jump_type448_wr              = ( waddr == JUMP_TYPE448_REG ) && wen;
wire jump_type449_wr              = ( waddr == JUMP_TYPE449_REG ) && wen;
wire jump_type450_wr              = ( waddr == JUMP_TYPE450_REG ) && wen;
wire jump_type451_wr              = ( waddr == JUMP_TYPE451_REG ) && wen;
wire jump_type452_wr              = ( waddr == JUMP_TYPE452_REG ) && wen;
wire jump_type453_wr              = ( waddr == JUMP_TYPE453_REG ) && wen;
wire jump_type454_wr              = ( waddr == JUMP_TYPE454_REG ) && wen;
wire jump_type455_wr              = ( waddr == JUMP_TYPE455_REG ) && wen;
wire jump_type456_wr              = ( waddr == JUMP_TYPE456_REG ) && wen;
wire jump_type457_wr              = ( waddr == JUMP_TYPE457_REG ) && wen;
wire jump_type458_wr              = ( waddr == JUMP_TYPE458_REG ) && wen;
wire jump_type459_wr              = ( waddr == JUMP_TYPE459_REG ) && wen;
wire jump_type460_wr              = ( waddr == JUMP_TYPE460_REG ) && wen;
wire jump_type461_wr              = ( waddr == JUMP_TYPE461_REG ) && wen;
wire jump_type462_wr              = ( waddr == JUMP_TYPE462_REG ) && wen;
wire jump_type463_wr              = ( waddr == JUMP_TYPE463_REG ) && wen;
wire jump_type464_wr              = ( waddr == JUMP_TYPE464_REG ) && wen;
wire jump_type465_wr              = ( waddr == JUMP_TYPE465_REG ) && wen;
wire jump_type466_wr              = ( waddr == JUMP_TYPE466_REG ) && wen;
wire jump_type467_wr              = ( waddr == JUMP_TYPE467_REG ) && wen;
wire jump_type468_wr              = ( waddr == JUMP_TYPE468_REG ) && wen;
wire jump_type469_wr              = ( waddr == JUMP_TYPE469_REG ) && wen;
wire jump_type470_wr              = ( waddr == JUMP_TYPE470_REG ) && wen;
wire jump_type471_wr              = ( waddr == JUMP_TYPE471_REG ) && wen;
wire jump_type472_wr              = ( waddr == JUMP_TYPE472_REG ) && wen;
wire jump_type473_wr              = ( waddr == JUMP_TYPE473_REG ) && wen;
wire jump_type474_wr              = ( waddr == JUMP_TYPE474_REG ) && wen;
wire jump_type475_wr              = ( waddr == JUMP_TYPE475_REG ) && wen;
wire jump_type476_wr              = ( waddr == JUMP_TYPE476_REG ) && wen;
wire jump_type477_wr              = ( waddr == JUMP_TYPE477_REG ) && wen;
wire jump_type478_wr              = ( waddr == JUMP_TYPE478_REG ) && wen;
wire jump_type479_wr              = ( waddr == JUMP_TYPE479_REG ) && wen;
wire jump_type480_wr              = ( waddr == JUMP_TYPE480_REG ) && wen;
wire jump_type481_wr              = ( waddr == JUMP_TYPE481_REG ) && wen;
wire jump_type482_wr              = ( waddr == JUMP_TYPE482_REG ) && wen;
wire jump_type483_wr              = ( waddr == JUMP_TYPE483_REG ) && wen;
wire jump_type484_wr              = ( waddr == JUMP_TYPE484_REG ) && wen;
wire jump_type485_wr              = ( waddr == JUMP_TYPE485_REG ) && wen;
wire jump_type486_wr              = ( waddr == JUMP_TYPE486_REG ) && wen;
wire jump_type487_wr              = ( waddr == JUMP_TYPE487_REG ) && wen;
wire jump_type488_wr              = ( waddr == JUMP_TYPE488_REG ) && wen;
wire jump_type489_wr              = ( waddr == JUMP_TYPE489_REG ) && wen;
wire jump_type490_wr              = ( waddr == JUMP_TYPE490_REG ) && wen;
wire jump_type491_wr              = ( waddr == JUMP_TYPE491_REG ) && wen;
wire jump_type492_wr              = ( waddr == JUMP_TYPE492_REG ) && wen;
wire jump_type493_wr              = ( waddr == JUMP_TYPE493_REG ) && wen;
wire jump_type494_wr              = ( waddr == JUMP_TYPE494_REG ) && wen;
wire jump_type495_wr              = ( waddr == JUMP_TYPE495_REG ) && wen;
wire jump_type496_wr              = ( waddr == JUMP_TYPE496_REG ) && wen;
wire jump_type497_wr              = ( waddr == JUMP_TYPE497_REG ) && wen;
wire jump_type498_wr              = ( waddr == JUMP_TYPE498_REG ) && wen;
wire jump_type499_wr              = ( waddr == JUMP_TYPE499_REG ) && wen;
wire jump_type500_wr              = ( waddr == JUMP_TYPE500_REG ) && wen;
wire jump_type501_wr              = ( waddr == JUMP_TYPE501_REG ) && wen;
wire jump_type502_wr              = ( waddr == JUMP_TYPE502_REG ) && wen;
wire jump_type503_wr              = ( waddr == JUMP_TYPE503_REG ) && wen;
wire jump_type504_wr              = ( waddr == JUMP_TYPE504_REG ) && wen;
wire jump_type505_wr              = ( waddr == JUMP_TYPE505_REG ) && wen;
wire jump_type506_wr              = ( waddr == JUMP_TYPE506_REG ) && wen;
wire jump_type507_wr              = ( waddr == JUMP_TYPE507_REG ) && wen;
wire jump_type508_wr              = ( waddr == JUMP_TYPE508_REG ) && wen;
wire jump_type509_wr              = ( waddr == JUMP_TYPE509_REG ) && wen;
wire jump_type510_wr              = ( waddr == JUMP_TYPE510_REG ) && wen;
wire jump_type511_wr              = ( waddr == JUMP_TYPE511_REG ) && wen;

//--------------------------------processing------------------------------------------------

//common_para
assign common_para_reg[31:26] = 6'h0                     ;
assign common_para_reg[25:24] = dcrc_num                 ;
assign common_para_reg[23:22] = list_num                 ;
assign common_para_reg[21]   = leaf_mode                ;
assign common_para_reg[20:12] = param_k                  ;
assign common_para_reg[11:3] = param_a                  ;
assign common_para_reg[2:0]  = param_n                  ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        dcrc_num <= 2'h0;
    else if( common_para_wr )
        dcrc_num <= wdata[25:24];
end

always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        list_num <= 2'h0;
    else if( common_para_wr )
        list_num <= wdata[23:22];
end

always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        leaf_mode <= 1'h0;
    else if( common_para_wr )
        leaf_mode <= wdata[21];
end

always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        param_k <= 9'h0;
    else if( common_para_wr )
        param_k <= wdata[20:12];
end

always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        param_a <= 9'h0;
    else if( common_para_wr )
        param_a <= wdata[11:3];
end

always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        param_n <= 3'h0;
    else if( common_para_wr )
        param_n <= wdata[2:0];
end


//jump_type0
assign jump_type0_reg[31:0]   = jump_type0                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type0 <= 32'h0;
    else if( jump_type0_wr )
        jump_type0 <= wdata[31:0];
end


//jump_type1
assign jump_type1_reg[31:0]   = jump_type1                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type1 <= 32'h0;
    else if( jump_type1_wr )
        jump_type1 <= wdata[31:0];
end


//jump_type2
assign jump_type2_reg[31:0]   = jump_type2                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type2 <= 32'h0;
    else if( jump_type2_wr )
        jump_type2 <= wdata[31:0];
end


//jump_type3
assign jump_type3_reg[31:0]   = jump_type3                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type3 <= 32'h0;
    else if( jump_type3_wr )
        jump_type3 <= wdata[31:0];
end


//jump_type4
assign jump_type4_reg[31:0]   = jump_type4                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type4 <= 32'h0;
    else if( jump_type4_wr )
        jump_type4 <= wdata[31:0];
end


//jump_type5
assign jump_type5_reg[31:0]   = jump_type5                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type5 <= 32'h0;
    else if( jump_type5_wr )
        jump_type5 <= wdata[31:0];
end


//jump_type6
assign jump_type6_reg[31:0]   = jump_type6                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type6 <= 32'h0;
    else if( jump_type6_wr )
        jump_type6 <= wdata[31:0];
end


//jump_type7
assign jump_type7_reg[31:0]   = jump_type7                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type7 <= 32'h0;
    else if( jump_type7_wr )
        jump_type7 <= wdata[31:0];
end


//jump_type8
assign jump_type8_reg[31:0]   = jump_type8                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type8 <= 32'h0;
    else if( jump_type8_wr )
        jump_type8 <= wdata[31:0];
end


//jump_type9
assign jump_type9_reg[31:0]   = jump_type9                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type9 <= 32'h0;
    else if( jump_type9_wr )
        jump_type9 <= wdata[31:0];
end


//jump_type10
assign jump_type10_reg[31:0]   = jump_type10                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type10 <= 32'h0;
    else if( jump_type10_wr )
        jump_type10 <= wdata[31:0];
end


//jump_type11
assign jump_type11_reg[31:0]   = jump_type11                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type11 <= 32'h0;
    else if( jump_type11_wr )
        jump_type11 <= wdata[31:0];
end


//jump_type12
assign jump_type12_reg[31:0]   = jump_type12                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type12 <= 32'h0;
    else if( jump_type12_wr )
        jump_type12 <= wdata[31:0];
end


//jump_type13
assign jump_type13_reg[31:0]   = jump_type13                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type13 <= 32'h0;
    else if( jump_type13_wr )
        jump_type13 <= wdata[31:0];
end


//jump_type14
assign jump_type14_reg[31:0]   = jump_type14                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type14 <= 32'h0;
    else if( jump_type14_wr )
        jump_type14 <= wdata[31:0];
end


//jump_type15
assign jump_type15_reg[31:0]   = jump_type15                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type15 <= 32'h0;
    else if( jump_type15_wr )
        jump_type15 <= wdata[31:0];
end


//jump_type16
assign jump_type16_reg[31:0]   = jump_type16                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type16 <= 32'h0;
    else if( jump_type16_wr )
        jump_type16 <= wdata[31:0];
end


//jump_type17
assign jump_type17_reg[31:0]   = jump_type17                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type17 <= 32'h0;
    else if( jump_type17_wr )
        jump_type17 <= wdata[31:0];
end


//jump_type18
assign jump_type18_reg[31:0]   = jump_type18                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type18 <= 32'h0;
    else if( jump_type18_wr )
        jump_type18 <= wdata[31:0];
end


//jump_type19
assign jump_type19_reg[31:0]   = jump_type19                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type19 <= 32'h0;
    else if( jump_type19_wr )
        jump_type19 <= wdata[31:0];
end


//jump_type20
assign jump_type20_reg[31:0]   = jump_type20                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type20 <= 32'h0;
    else if( jump_type20_wr )
        jump_type20 <= wdata[31:0];
end


//jump_type21
assign jump_type21_reg[31:0]   = jump_type21                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type21 <= 32'h0;
    else if( jump_type21_wr )
        jump_type21 <= wdata[31:0];
end


//jump_type22
assign jump_type22_reg[31:0]   = jump_type22                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type22 <= 32'h0;
    else if( jump_type22_wr )
        jump_type22 <= wdata[31:0];
end


//jump_type23
assign jump_type23_reg[31:0]   = jump_type23                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type23 <= 32'h0;
    else if( jump_type23_wr )
        jump_type23 <= wdata[31:0];
end


//jump_type24
assign jump_type24_reg[31:0]   = jump_type24                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type24 <= 32'h0;
    else if( jump_type24_wr )
        jump_type24 <= wdata[31:0];
end


//jump_type25
assign jump_type25_reg[31:0]   = jump_type25                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type25 <= 32'h0;
    else if( jump_type25_wr )
        jump_type25 <= wdata[31:0];
end


//jump_type26
assign jump_type26_reg[31:0]   = jump_type26                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type26 <= 32'h0;
    else if( jump_type26_wr )
        jump_type26 <= wdata[31:0];
end


//jump_type27
assign jump_type27_reg[31:0]   = jump_type27                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type27 <= 32'h0;
    else if( jump_type27_wr )
        jump_type27 <= wdata[31:0];
end


//jump_type28
assign jump_type28_reg[31:0]   = jump_type28                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type28 <= 32'h0;
    else if( jump_type28_wr )
        jump_type28 <= wdata[31:0];
end


//jump_type29
assign jump_type29_reg[31:0]   = jump_type29                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type29 <= 32'h0;
    else if( jump_type29_wr )
        jump_type29 <= wdata[31:0];
end


//jump_type30
assign jump_type30_reg[31:0]   = jump_type30                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type30 <= 32'h0;
    else if( jump_type30_wr )
        jump_type30 <= wdata[31:0];
end


//jump_type31
assign jump_type31_reg[31:0]   = jump_type31                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type31 <= 32'h0;
    else if( jump_type31_wr )
        jump_type31 <= wdata[31:0];
end


//jump_type32
assign jump_type32_reg[31:0]   = jump_type32                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type32 <= 32'h0;
    else if( jump_type32_wr )
        jump_type32 <= wdata[31:0];
end


//jump_type33
assign jump_type33_reg[31:0]   = jump_type33                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type33 <= 32'h0;
    else if( jump_type33_wr )
        jump_type33 <= wdata[31:0];
end


//jump_type34
assign jump_type34_reg[31:0]   = jump_type34                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type34 <= 32'h0;
    else if( jump_type34_wr )
        jump_type34 <= wdata[31:0];
end


//jump_type35
assign jump_type35_reg[31:0]   = jump_type35                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type35 <= 32'h0;
    else if( jump_type35_wr )
        jump_type35 <= wdata[31:0];
end


//jump_type36
assign jump_type36_reg[31:0]   = jump_type36                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type36 <= 32'h0;
    else if( jump_type36_wr )
        jump_type36 <= wdata[31:0];
end


//jump_type37
assign jump_type37_reg[31:0]   = jump_type37                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type37 <= 32'h0;
    else if( jump_type37_wr )
        jump_type37 <= wdata[31:0];
end


//jump_type38
assign jump_type38_reg[31:0]   = jump_type38                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type38 <= 32'h0;
    else if( jump_type38_wr )
        jump_type38 <= wdata[31:0];
end


//jump_type39
assign jump_type39_reg[31:0]   = jump_type39                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type39 <= 32'h0;
    else if( jump_type39_wr )
        jump_type39 <= wdata[31:0];
end


//jump_type40
assign jump_type40_reg[31:0]   = jump_type40                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type40 <= 32'h0;
    else if( jump_type40_wr )
        jump_type40 <= wdata[31:0];
end


//jump_type41
assign jump_type41_reg[31:0]   = jump_type41                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type41 <= 32'h0;
    else if( jump_type41_wr )
        jump_type41 <= wdata[31:0];
end


//jump_type42
assign jump_type42_reg[31:0]   = jump_type42                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type42 <= 32'h0;
    else if( jump_type42_wr )
        jump_type42 <= wdata[31:0];
end


//jump_type43
assign jump_type43_reg[31:0]   = jump_type43                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type43 <= 32'h0;
    else if( jump_type43_wr )
        jump_type43 <= wdata[31:0];
end


//jump_type44
assign jump_type44_reg[31:0]   = jump_type44                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type44 <= 32'h0;
    else if( jump_type44_wr )
        jump_type44 <= wdata[31:0];
end


//jump_type45
assign jump_type45_reg[31:0]   = jump_type45                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type45 <= 32'h0;
    else if( jump_type45_wr )
        jump_type45 <= wdata[31:0];
end


//jump_type46
assign jump_type46_reg[31:0]   = jump_type46                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type46 <= 32'h0;
    else if( jump_type46_wr )
        jump_type46 <= wdata[31:0];
end


//jump_type47
assign jump_type47_reg[31:0]   = jump_type47                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type47 <= 32'h0;
    else if( jump_type47_wr )
        jump_type47 <= wdata[31:0];
end


//jump_type48
assign jump_type48_reg[31:0]   = jump_type48                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type48 <= 32'h0;
    else if( jump_type48_wr )
        jump_type48 <= wdata[31:0];
end


//jump_type49
assign jump_type49_reg[31:0]   = jump_type49                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type49 <= 32'h0;
    else if( jump_type49_wr )
        jump_type49 <= wdata[31:0];
end


//jump_type50
assign jump_type50_reg[31:0]   = jump_type50                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type50 <= 32'h0;
    else if( jump_type50_wr )
        jump_type50 <= wdata[31:0];
end


//jump_type51
assign jump_type51_reg[31:0]   = jump_type51                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type51 <= 32'h0;
    else if( jump_type51_wr )
        jump_type51 <= wdata[31:0];
end


//jump_type52
assign jump_type52_reg[31:0]   = jump_type52                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type52 <= 32'h0;
    else if( jump_type52_wr )
        jump_type52 <= wdata[31:0];
end


//jump_type53
assign jump_type53_reg[31:0]   = jump_type53                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type53 <= 32'h0;
    else if( jump_type53_wr )
        jump_type53 <= wdata[31:0];
end


//jump_type54
assign jump_type54_reg[31:0]   = jump_type54                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type54 <= 32'h0;
    else if( jump_type54_wr )
        jump_type54 <= wdata[31:0];
end


//jump_type55
assign jump_type55_reg[31:0]   = jump_type55                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type55 <= 32'h0;
    else if( jump_type55_wr )
        jump_type55 <= wdata[31:0];
end


//jump_type56
assign jump_type56_reg[31:0]   = jump_type56                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type56 <= 32'h0;
    else if( jump_type56_wr )
        jump_type56 <= wdata[31:0];
end


//jump_type57
assign jump_type57_reg[31:0]   = jump_type57                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type57 <= 32'h0;
    else if( jump_type57_wr )
        jump_type57 <= wdata[31:0];
end


//jump_type58
assign jump_type58_reg[31:0]   = jump_type58                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type58 <= 32'h0;
    else if( jump_type58_wr )
        jump_type58 <= wdata[31:0];
end


//jump_type59
assign jump_type59_reg[31:0]   = jump_type59                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type59 <= 32'h0;
    else if( jump_type59_wr )
        jump_type59 <= wdata[31:0];
end


//jump_type60
assign jump_type60_reg[31:0]   = jump_type60                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type60 <= 32'h0;
    else if( jump_type60_wr )
        jump_type60 <= wdata[31:0];
end


//jump_type61
assign jump_type61_reg[31:0]   = jump_type61                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type61 <= 32'h0;
    else if( jump_type61_wr )
        jump_type61 <= wdata[31:0];
end


//jump_type62
assign jump_type62_reg[31:0]   = jump_type62                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type62 <= 32'h0;
    else if( jump_type62_wr )
        jump_type62 <= wdata[31:0];
end


//jump_type63
assign jump_type63_reg[31:0]   = jump_type63                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type63 <= 32'h0;
    else if( jump_type63_wr )
        jump_type63 <= wdata[31:0];
end


//jump_type64
assign jump_type64_reg[31:0]   = jump_type64                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type64 <= 32'h0;
    else if( jump_type64_wr )
        jump_type64 <= wdata[31:0];
end


//jump_type65
assign jump_type65_reg[31:0]   = jump_type65                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type65 <= 32'h0;
    else if( jump_type65_wr )
        jump_type65 <= wdata[31:0];
end


//jump_type66
assign jump_type66_reg[31:0]   = jump_type66                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type66 <= 32'h0;
    else if( jump_type66_wr )
        jump_type66 <= wdata[31:0];
end


//jump_type67
assign jump_type67_reg[31:0]   = jump_type67                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type67 <= 32'h0;
    else if( jump_type67_wr )
        jump_type67 <= wdata[31:0];
end


//jump_type68
assign jump_type68_reg[31:0]   = jump_type68                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type68 <= 32'h0;
    else if( jump_type68_wr )
        jump_type68 <= wdata[31:0];
end


//jump_type69
assign jump_type69_reg[31:0]   = jump_type69                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type69 <= 32'h0;
    else if( jump_type69_wr )
        jump_type69 <= wdata[31:0];
end


//jump_type70
assign jump_type70_reg[31:0]   = jump_type70                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type70 <= 32'h0;
    else if( jump_type70_wr )
        jump_type70 <= wdata[31:0];
end


//jump_type71
assign jump_type71_reg[31:0]   = jump_type71                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type71 <= 32'h0;
    else if( jump_type71_wr )
        jump_type71 <= wdata[31:0];
end


//jump_type72
assign jump_type72_reg[31:0]   = jump_type72                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type72 <= 32'h0;
    else if( jump_type72_wr )
        jump_type72 <= wdata[31:0];
end


//jump_type73
assign jump_type73_reg[31:0]   = jump_type73                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type73 <= 32'h0;
    else if( jump_type73_wr )
        jump_type73 <= wdata[31:0];
end


//jump_type74
assign jump_type74_reg[31:0]   = jump_type74                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type74 <= 32'h0;
    else if( jump_type74_wr )
        jump_type74 <= wdata[31:0];
end


//jump_type75
assign jump_type75_reg[31:0]   = jump_type75                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type75 <= 32'h0;
    else if( jump_type75_wr )
        jump_type75 <= wdata[31:0];
end


//jump_type76
assign jump_type76_reg[31:0]   = jump_type76                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type76 <= 32'h0;
    else if( jump_type76_wr )
        jump_type76 <= wdata[31:0];
end


//jump_type77
assign jump_type77_reg[31:0]   = jump_type77                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type77 <= 32'h0;
    else if( jump_type77_wr )
        jump_type77 <= wdata[31:0];
end


//jump_type78
assign jump_type78_reg[31:0]   = jump_type78                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type78 <= 32'h0;
    else if( jump_type78_wr )
        jump_type78 <= wdata[31:0];
end


//jump_type79
assign jump_type79_reg[31:0]   = jump_type79                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type79 <= 32'h0;
    else if( jump_type79_wr )
        jump_type79 <= wdata[31:0];
end


//jump_type80
assign jump_type80_reg[31:0]   = jump_type80                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type80 <= 32'h0;
    else if( jump_type80_wr )
        jump_type80 <= wdata[31:0];
end


//jump_type81
assign jump_type81_reg[31:0]   = jump_type81                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type81 <= 32'h0;
    else if( jump_type81_wr )
        jump_type81 <= wdata[31:0];
end


//jump_type82
assign jump_type82_reg[31:0]   = jump_type82                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type82 <= 32'h0;
    else if( jump_type82_wr )
        jump_type82 <= wdata[31:0];
end


//jump_type83
assign jump_type83_reg[31:0]   = jump_type83                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type83 <= 32'h0;
    else if( jump_type83_wr )
        jump_type83 <= wdata[31:0];
end


//jump_type84
assign jump_type84_reg[31:0]   = jump_type84                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type84 <= 32'h0;
    else if( jump_type84_wr )
        jump_type84 <= wdata[31:0];
end


//jump_type85
assign jump_type85_reg[31:0]   = jump_type85                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type85 <= 32'h0;
    else if( jump_type85_wr )
        jump_type85 <= wdata[31:0];
end


//jump_type86
assign jump_type86_reg[31:0]   = jump_type86                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type86 <= 32'h0;
    else if( jump_type86_wr )
        jump_type86 <= wdata[31:0];
end


//jump_type87
assign jump_type87_reg[31:0]   = jump_type87                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type87 <= 32'h0;
    else if( jump_type87_wr )
        jump_type87 <= wdata[31:0];
end


//jump_type88
assign jump_type88_reg[31:0]   = jump_type88                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type88 <= 32'h0;
    else if( jump_type88_wr )
        jump_type88 <= wdata[31:0];
end


//jump_type89
assign jump_type89_reg[31:0]   = jump_type89                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type89 <= 32'h0;
    else if( jump_type89_wr )
        jump_type89 <= wdata[31:0];
end


//jump_type90
assign jump_type90_reg[31:0]   = jump_type90                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type90 <= 32'h0;
    else if( jump_type90_wr )
        jump_type90 <= wdata[31:0];
end


//jump_type91
assign jump_type91_reg[31:0]   = jump_type91                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type91 <= 32'h0;
    else if( jump_type91_wr )
        jump_type91 <= wdata[31:0];
end


//jump_type92
assign jump_type92_reg[31:0]   = jump_type92                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type92 <= 32'h0;
    else if( jump_type92_wr )
        jump_type92 <= wdata[31:0];
end


//jump_type93
assign jump_type93_reg[31:0]   = jump_type93                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type93 <= 32'h0;
    else if( jump_type93_wr )
        jump_type93 <= wdata[31:0];
end


//jump_type94
assign jump_type94_reg[31:0]   = jump_type94                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type94 <= 32'h0;
    else if( jump_type94_wr )
        jump_type94 <= wdata[31:0];
end


//jump_type95
assign jump_type95_reg[31:0]   = jump_type95                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type95 <= 32'h0;
    else if( jump_type95_wr )
        jump_type95 <= wdata[31:0];
end


//jump_type96
assign jump_type96_reg[31:0]   = jump_type96                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type96 <= 32'h0;
    else if( jump_type96_wr )
        jump_type96 <= wdata[31:0];
end


//jump_type97
assign jump_type97_reg[31:0]   = jump_type97                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type97 <= 32'h0;
    else if( jump_type97_wr )
        jump_type97 <= wdata[31:0];
end


//jump_type98
assign jump_type98_reg[31:0]   = jump_type98                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type98 <= 32'h0;
    else if( jump_type98_wr )
        jump_type98 <= wdata[31:0];
end


//jump_type99
assign jump_type99_reg[31:0]   = jump_type99                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type99 <= 32'h0;
    else if( jump_type99_wr )
        jump_type99 <= wdata[31:0];
end


//jump_type100
assign jump_type100_reg[31:0]   = jump_type100                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type100 <= 32'h0;
    else if( jump_type100_wr )
        jump_type100 <= wdata[31:0];
end


//jump_type101
assign jump_type101_reg[31:0]   = jump_type101                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type101 <= 32'h0;
    else if( jump_type101_wr )
        jump_type101 <= wdata[31:0];
end


//jump_type102
assign jump_type102_reg[31:0]   = jump_type102                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type102 <= 32'h0;
    else if( jump_type102_wr )
        jump_type102 <= wdata[31:0];
end


//jump_type103
assign jump_type103_reg[31:0]   = jump_type103                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type103 <= 32'h0;
    else if( jump_type103_wr )
        jump_type103 <= wdata[31:0];
end


//jump_type104
assign jump_type104_reg[31:0]   = jump_type104                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type104 <= 32'h0;
    else if( jump_type104_wr )
        jump_type104 <= wdata[31:0];
end


//jump_type105
assign jump_type105_reg[31:0]   = jump_type105                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type105 <= 32'h0;
    else if( jump_type105_wr )
        jump_type105 <= wdata[31:0];
end


//jump_type106
assign jump_type106_reg[31:0]   = jump_type106                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type106 <= 32'h0;
    else if( jump_type106_wr )
        jump_type106 <= wdata[31:0];
end


//jump_type107
assign jump_type107_reg[31:0]   = jump_type107                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type107 <= 32'h0;
    else if( jump_type107_wr )
        jump_type107 <= wdata[31:0];
end


//jump_type108
assign jump_type108_reg[31:0]   = jump_type108                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type108 <= 32'h0;
    else if( jump_type108_wr )
        jump_type108 <= wdata[31:0];
end


//jump_type109
assign jump_type109_reg[31:0]   = jump_type109                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type109 <= 32'h0;
    else if( jump_type109_wr )
        jump_type109 <= wdata[31:0];
end


//jump_type110
assign jump_type110_reg[31:0]   = jump_type110                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type110 <= 32'h0;
    else if( jump_type110_wr )
        jump_type110 <= wdata[31:0];
end


//jump_type111
assign jump_type111_reg[31:0]   = jump_type111                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type111 <= 32'h0;
    else if( jump_type111_wr )
        jump_type111 <= wdata[31:0];
end


//jump_type112
assign jump_type112_reg[31:0]   = jump_type112                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type112 <= 32'h0;
    else if( jump_type112_wr )
        jump_type112 <= wdata[31:0];
end


//jump_type113
assign jump_type113_reg[31:0]   = jump_type113                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type113 <= 32'h0;
    else if( jump_type113_wr )
        jump_type113 <= wdata[31:0];
end


//jump_type114
assign jump_type114_reg[31:0]   = jump_type114                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type114 <= 32'h0;
    else if( jump_type114_wr )
        jump_type114 <= wdata[31:0];
end


//jump_type115
assign jump_type115_reg[31:0]   = jump_type115                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type115 <= 32'h0;
    else if( jump_type115_wr )
        jump_type115 <= wdata[31:0];
end


//jump_type116
assign jump_type116_reg[31:0]   = jump_type116                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type116 <= 32'h0;
    else if( jump_type116_wr )
        jump_type116 <= wdata[31:0];
end


//jump_type117
assign jump_type117_reg[31:0]   = jump_type117                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type117 <= 32'h0;
    else if( jump_type117_wr )
        jump_type117 <= wdata[31:0];
end


//jump_type118
assign jump_type118_reg[31:0]   = jump_type118                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type118 <= 32'h0;
    else if( jump_type118_wr )
        jump_type118 <= wdata[31:0];
end


//jump_type119
assign jump_type119_reg[31:0]   = jump_type119                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type119 <= 32'h0;
    else if( jump_type119_wr )
        jump_type119 <= wdata[31:0];
end


//jump_type120
assign jump_type120_reg[31:0]   = jump_type120                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type120 <= 32'h0;
    else if( jump_type120_wr )
        jump_type120 <= wdata[31:0];
end


//jump_type121
assign jump_type121_reg[31:0]   = jump_type121                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type121 <= 32'h0;
    else if( jump_type121_wr )
        jump_type121 <= wdata[31:0];
end


//jump_type122
assign jump_type122_reg[31:0]   = jump_type122                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type122 <= 32'h0;
    else if( jump_type122_wr )
        jump_type122 <= wdata[31:0];
end


//jump_type123
assign jump_type123_reg[31:0]   = jump_type123                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type123 <= 32'h0;
    else if( jump_type123_wr )
        jump_type123 <= wdata[31:0];
end


//jump_type124
assign jump_type124_reg[31:0]   = jump_type124                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type124 <= 32'h0;
    else if( jump_type124_wr )
        jump_type124 <= wdata[31:0];
end


//jump_type125
assign jump_type125_reg[31:0]   = jump_type125                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type125 <= 32'h0;
    else if( jump_type125_wr )
        jump_type125 <= wdata[31:0];
end


//jump_type126
assign jump_type126_reg[31:0]   = jump_type126                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type126 <= 32'h0;
    else if( jump_type126_wr )
        jump_type126 <= wdata[31:0];
end


//jump_type127
assign jump_type127_reg[31:0]   = jump_type127                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type127 <= 32'h0;
    else if( jump_type127_wr )
        jump_type127 <= wdata[31:0];
end


//jump_type128
assign jump_type128_reg[31:0]   = jump_type128                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type128 <= 32'h0;
    else if( jump_type128_wr )
        jump_type128 <= wdata[31:0];
end


//jump_type129
assign jump_type129_reg[31:0]   = jump_type129                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type129 <= 32'h0;
    else if( jump_type129_wr )
        jump_type129 <= wdata[31:0];
end


//jump_type130
assign jump_type130_reg[31:0]   = jump_type130                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type130 <= 32'h0;
    else if( jump_type130_wr )
        jump_type130 <= wdata[31:0];
end


//jump_type131
assign jump_type131_reg[31:0]   = jump_type131                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type131 <= 32'h0;
    else if( jump_type131_wr )
        jump_type131 <= wdata[31:0];
end


//jump_type132
assign jump_type132_reg[31:0]   = jump_type132                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type132 <= 32'h0;
    else if( jump_type132_wr )
        jump_type132 <= wdata[31:0];
end


//jump_type133
assign jump_type133_reg[31:0]   = jump_type133                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type133 <= 32'h0;
    else if( jump_type133_wr )
        jump_type133 <= wdata[31:0];
end


//jump_type134
assign jump_type134_reg[31:0]   = jump_type134                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type134 <= 32'h0;
    else if( jump_type134_wr )
        jump_type134 <= wdata[31:0];
end


//jump_type135
assign jump_type135_reg[31:0]   = jump_type135                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type135 <= 32'h0;
    else if( jump_type135_wr )
        jump_type135 <= wdata[31:0];
end


//jump_type136
assign jump_type136_reg[31:0]   = jump_type136                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type136 <= 32'h0;
    else if( jump_type136_wr )
        jump_type136 <= wdata[31:0];
end


//jump_type137
assign jump_type137_reg[31:0]   = jump_type137                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type137 <= 32'h0;
    else if( jump_type137_wr )
        jump_type137 <= wdata[31:0];
end


//jump_type138
assign jump_type138_reg[31:0]   = jump_type138                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type138 <= 32'h0;
    else if( jump_type138_wr )
        jump_type138 <= wdata[31:0];
end


//jump_type139
assign jump_type139_reg[31:0]   = jump_type139                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type139 <= 32'h0;
    else if( jump_type139_wr )
        jump_type139 <= wdata[31:0];
end


//jump_type140
assign jump_type140_reg[31:0]   = jump_type140                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type140 <= 32'h0;
    else if( jump_type140_wr )
        jump_type140 <= wdata[31:0];
end


//jump_type141
assign jump_type141_reg[31:0]   = jump_type141                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type141 <= 32'h0;
    else if( jump_type141_wr )
        jump_type141 <= wdata[31:0];
end


//jump_type142
assign jump_type142_reg[31:0]   = jump_type142                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type142 <= 32'h0;
    else if( jump_type142_wr )
        jump_type142 <= wdata[31:0];
end


//jump_type143
assign jump_type143_reg[31:0]   = jump_type143                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type143 <= 32'h0;
    else if( jump_type143_wr )
        jump_type143 <= wdata[31:0];
end


//jump_type144
assign jump_type144_reg[31:0]   = jump_type144                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type144 <= 32'h0;
    else if( jump_type144_wr )
        jump_type144 <= wdata[31:0];
end


//jump_type145
assign jump_type145_reg[31:0]   = jump_type145                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type145 <= 32'h0;
    else if( jump_type145_wr )
        jump_type145 <= wdata[31:0];
end


//jump_type146
assign jump_type146_reg[31:0]   = jump_type146                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type146 <= 32'h0;
    else if( jump_type146_wr )
        jump_type146 <= wdata[31:0];
end


//jump_type147
assign jump_type147_reg[31:0]   = jump_type147                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type147 <= 32'h0;
    else if( jump_type147_wr )
        jump_type147 <= wdata[31:0];
end


//jump_type148
assign jump_type148_reg[31:0]   = jump_type148                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type148 <= 32'h0;
    else if( jump_type148_wr )
        jump_type148 <= wdata[31:0];
end


//jump_type149
assign jump_type149_reg[31:0]   = jump_type149                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type149 <= 32'h0;
    else if( jump_type149_wr )
        jump_type149 <= wdata[31:0];
end


//jump_type150
assign jump_type150_reg[31:0]   = jump_type150                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type150 <= 32'h0;
    else if( jump_type150_wr )
        jump_type150 <= wdata[31:0];
end


//jump_type151
assign jump_type151_reg[31:0]   = jump_type151                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type151 <= 32'h0;
    else if( jump_type151_wr )
        jump_type151 <= wdata[31:0];
end


//jump_type152
assign jump_type152_reg[31:0]   = jump_type152                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type152 <= 32'h0;
    else if( jump_type152_wr )
        jump_type152 <= wdata[31:0];
end


//jump_type153
assign jump_type153_reg[31:0]   = jump_type153                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type153 <= 32'h0;
    else if( jump_type153_wr )
        jump_type153 <= wdata[31:0];
end


//jump_type154
assign jump_type154_reg[31:0]   = jump_type154                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type154 <= 32'h0;
    else if( jump_type154_wr )
        jump_type154 <= wdata[31:0];
end


//jump_type155
assign jump_type155_reg[31:0]   = jump_type155                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type155 <= 32'h0;
    else if( jump_type155_wr )
        jump_type155 <= wdata[31:0];
end


//jump_type156
assign jump_type156_reg[31:0]   = jump_type156                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type156 <= 32'h0;
    else if( jump_type156_wr )
        jump_type156 <= wdata[31:0];
end


//jump_type157
assign jump_type157_reg[31:0]   = jump_type157                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type157 <= 32'h0;
    else if( jump_type157_wr )
        jump_type157 <= wdata[31:0];
end


//jump_type158
assign jump_type158_reg[31:0]   = jump_type158                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type158 <= 32'h0;
    else if( jump_type158_wr )
        jump_type158 <= wdata[31:0];
end


//jump_type159
assign jump_type159_reg[31:0]   = jump_type159                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type159 <= 32'h0;
    else if( jump_type159_wr )
        jump_type159 <= wdata[31:0];
end


//jump_type160
assign jump_type160_reg[31:0]   = jump_type160                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type160 <= 32'h0;
    else if( jump_type160_wr )
        jump_type160 <= wdata[31:0];
end


//jump_type161
assign jump_type161_reg[31:0]   = jump_type161                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type161 <= 32'h0;
    else if( jump_type161_wr )
        jump_type161 <= wdata[31:0];
end


//jump_type162
assign jump_type162_reg[31:0]   = jump_type162                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type162 <= 32'h0;
    else if( jump_type162_wr )
        jump_type162 <= wdata[31:0];
end


//jump_type163
assign jump_type163_reg[31:0]   = jump_type163                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type163 <= 32'h0;
    else if( jump_type163_wr )
        jump_type163 <= wdata[31:0];
end


//jump_type164
assign jump_type164_reg[31:0]   = jump_type164                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type164 <= 32'h0;
    else if( jump_type164_wr )
        jump_type164 <= wdata[31:0];
end


//jump_type165
assign jump_type165_reg[31:0]   = jump_type165                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type165 <= 32'h0;
    else if( jump_type165_wr )
        jump_type165 <= wdata[31:0];
end


//jump_type166
assign jump_type166_reg[31:0]   = jump_type166                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type166 <= 32'h0;
    else if( jump_type166_wr )
        jump_type166 <= wdata[31:0];
end


//jump_type167
assign jump_type167_reg[31:0]   = jump_type167                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type167 <= 32'h0;
    else if( jump_type167_wr )
        jump_type167 <= wdata[31:0];
end


//jump_type168
assign jump_type168_reg[31:0]   = jump_type168                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type168 <= 32'h0;
    else if( jump_type168_wr )
        jump_type168 <= wdata[31:0];
end


//jump_type169
assign jump_type169_reg[31:0]   = jump_type169                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type169 <= 32'h0;
    else if( jump_type169_wr )
        jump_type169 <= wdata[31:0];
end


//jump_type170
assign jump_type170_reg[31:0]   = jump_type170                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type170 <= 32'h0;
    else if( jump_type170_wr )
        jump_type170 <= wdata[31:0];
end


//jump_type171
assign jump_type171_reg[31:0]   = jump_type171                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type171 <= 32'h0;
    else if( jump_type171_wr )
        jump_type171 <= wdata[31:0];
end


//jump_type172
assign jump_type172_reg[31:0]   = jump_type172                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type172 <= 32'h0;
    else if( jump_type172_wr )
        jump_type172 <= wdata[31:0];
end


//jump_type173
assign jump_type173_reg[31:0]   = jump_type173                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type173 <= 32'h0;
    else if( jump_type173_wr )
        jump_type173 <= wdata[31:0];
end


//jump_type174
assign jump_type174_reg[31:0]   = jump_type174                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type174 <= 32'h0;
    else if( jump_type174_wr )
        jump_type174 <= wdata[31:0];
end


//jump_type175
assign jump_type175_reg[31:0]   = jump_type175                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type175 <= 32'h0;
    else if( jump_type175_wr )
        jump_type175 <= wdata[31:0];
end


//jump_type176
assign jump_type176_reg[31:0]   = jump_type176                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type176 <= 32'h0;
    else if( jump_type176_wr )
        jump_type176 <= wdata[31:0];
end


//jump_type177
assign jump_type177_reg[31:0]   = jump_type177                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type177 <= 32'h0;
    else if( jump_type177_wr )
        jump_type177 <= wdata[31:0];
end


//jump_type178
assign jump_type178_reg[31:0]   = jump_type178                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type178 <= 32'h0;
    else if( jump_type178_wr )
        jump_type178 <= wdata[31:0];
end


//jump_type179
assign jump_type179_reg[31:0]   = jump_type179                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type179 <= 32'h0;
    else if( jump_type179_wr )
        jump_type179 <= wdata[31:0];
end


//jump_type180
assign jump_type180_reg[31:0]   = jump_type180                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type180 <= 32'h0;
    else if( jump_type180_wr )
        jump_type180 <= wdata[31:0];
end


//jump_type181
assign jump_type181_reg[31:0]   = jump_type181                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type181 <= 32'h0;
    else if( jump_type181_wr )
        jump_type181 <= wdata[31:0];
end


//jump_type182
assign jump_type182_reg[31:0]   = jump_type182                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type182 <= 32'h0;
    else if( jump_type182_wr )
        jump_type182 <= wdata[31:0];
end


//jump_type183
assign jump_type183_reg[31:0]   = jump_type183                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type183 <= 32'h0;
    else if( jump_type183_wr )
        jump_type183 <= wdata[31:0];
end


//jump_type184
assign jump_type184_reg[31:0]   = jump_type184                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type184 <= 32'h0;
    else if( jump_type184_wr )
        jump_type184 <= wdata[31:0];
end


//jump_type185
assign jump_type185_reg[31:0]   = jump_type185                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type185 <= 32'h0;
    else if( jump_type185_wr )
        jump_type185 <= wdata[31:0];
end


//jump_type186
assign jump_type186_reg[31:0]   = jump_type186                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type186 <= 32'h0;
    else if( jump_type186_wr )
        jump_type186 <= wdata[31:0];
end


//jump_type187
assign jump_type187_reg[31:0]   = jump_type187                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type187 <= 32'h0;
    else if( jump_type187_wr )
        jump_type187 <= wdata[31:0];
end


//jump_type188
assign jump_type188_reg[31:0]   = jump_type188                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type188 <= 32'h0;
    else if( jump_type188_wr )
        jump_type188 <= wdata[31:0];
end


//jump_type189
assign jump_type189_reg[31:0]   = jump_type189                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type189 <= 32'h0;
    else if( jump_type189_wr )
        jump_type189 <= wdata[31:0];
end


//jump_type190
assign jump_type190_reg[31:0]   = jump_type190                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type190 <= 32'h0;
    else if( jump_type190_wr )
        jump_type190 <= wdata[31:0];
end


//jump_type191
assign jump_type191_reg[31:0]   = jump_type191                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type191 <= 32'h0;
    else if( jump_type191_wr )
        jump_type191 <= wdata[31:0];
end


//jump_type192
assign jump_type192_reg[31:0]   = jump_type192                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type192 <= 32'h0;
    else if( jump_type192_wr )
        jump_type192 <= wdata[31:0];
end


//jump_type193
assign jump_type193_reg[31:0]   = jump_type193                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type193 <= 32'h0;
    else if( jump_type193_wr )
        jump_type193 <= wdata[31:0];
end


//jump_type194
assign jump_type194_reg[31:0]   = jump_type194                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type194 <= 32'h0;
    else if( jump_type194_wr )
        jump_type194 <= wdata[31:0];
end


//jump_type195
assign jump_type195_reg[31:0]   = jump_type195                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type195 <= 32'h0;
    else if( jump_type195_wr )
        jump_type195 <= wdata[31:0];
end


//jump_type196
assign jump_type196_reg[31:0]   = jump_type196                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type196 <= 32'h0;
    else if( jump_type196_wr )
        jump_type196 <= wdata[31:0];
end


//jump_type197
assign jump_type197_reg[31:0]   = jump_type197                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type197 <= 32'h0;
    else if( jump_type197_wr )
        jump_type197 <= wdata[31:0];
end


//jump_type198
assign jump_type198_reg[31:0]   = jump_type198                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type198 <= 32'h0;
    else if( jump_type198_wr )
        jump_type198 <= wdata[31:0];
end


//jump_type199
assign jump_type199_reg[31:0]   = jump_type199                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type199 <= 32'h0;
    else if( jump_type199_wr )
        jump_type199 <= wdata[31:0];
end


//jump_type200
assign jump_type200_reg[31:0]   = jump_type200                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type200 <= 32'h0;
    else if( jump_type200_wr )
        jump_type200 <= wdata[31:0];
end


//jump_type201
assign jump_type201_reg[31:0]   = jump_type201                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type201 <= 32'h0;
    else if( jump_type201_wr )
        jump_type201 <= wdata[31:0];
end


//jump_type202
assign jump_type202_reg[31:0]   = jump_type202                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type202 <= 32'h0;
    else if( jump_type202_wr )
        jump_type202 <= wdata[31:0];
end


//jump_type203
assign jump_type203_reg[31:0]   = jump_type203                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type203 <= 32'h0;
    else if( jump_type203_wr )
        jump_type203 <= wdata[31:0];
end


//jump_type204
assign jump_type204_reg[31:0]   = jump_type204                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type204 <= 32'h0;
    else if( jump_type204_wr )
        jump_type204 <= wdata[31:0];
end


//jump_type205
assign jump_type205_reg[31:0]   = jump_type205                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type205 <= 32'h0;
    else if( jump_type205_wr )
        jump_type205 <= wdata[31:0];
end


//jump_type206
assign jump_type206_reg[31:0]   = jump_type206                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type206 <= 32'h0;
    else if( jump_type206_wr )
        jump_type206 <= wdata[31:0];
end


//jump_type207
assign jump_type207_reg[31:0]   = jump_type207                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type207 <= 32'h0;
    else if( jump_type207_wr )
        jump_type207 <= wdata[31:0];
end


//jump_type208
assign jump_type208_reg[31:0]   = jump_type208                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type208 <= 32'h0;
    else if( jump_type208_wr )
        jump_type208 <= wdata[31:0];
end


//jump_type209
assign jump_type209_reg[31:0]   = jump_type209                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type209 <= 32'h0;
    else if( jump_type209_wr )
        jump_type209 <= wdata[31:0];
end


//jump_type210
assign jump_type210_reg[31:0]   = jump_type210                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type210 <= 32'h0;
    else if( jump_type210_wr )
        jump_type210 <= wdata[31:0];
end


//jump_type211
assign jump_type211_reg[31:0]   = jump_type211                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type211 <= 32'h0;
    else if( jump_type211_wr )
        jump_type211 <= wdata[31:0];
end


//jump_type212
assign jump_type212_reg[31:0]   = jump_type212                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type212 <= 32'h0;
    else if( jump_type212_wr )
        jump_type212 <= wdata[31:0];
end


//jump_type213
assign jump_type213_reg[31:0]   = jump_type213                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type213 <= 32'h0;
    else if( jump_type213_wr )
        jump_type213 <= wdata[31:0];
end


//jump_type214
assign jump_type214_reg[31:0]   = jump_type214                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type214 <= 32'h0;
    else if( jump_type214_wr )
        jump_type214 <= wdata[31:0];
end


//jump_type215
assign jump_type215_reg[31:0]   = jump_type215                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type215 <= 32'h0;
    else if( jump_type215_wr )
        jump_type215 <= wdata[31:0];
end


//jump_type216
assign jump_type216_reg[31:0]   = jump_type216                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type216 <= 32'h0;
    else if( jump_type216_wr )
        jump_type216 <= wdata[31:0];
end


//jump_type217
assign jump_type217_reg[31:0]   = jump_type217                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type217 <= 32'h0;
    else if( jump_type217_wr )
        jump_type217 <= wdata[31:0];
end


//jump_type218
assign jump_type218_reg[31:0]   = jump_type218                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type218 <= 32'h0;
    else if( jump_type218_wr )
        jump_type218 <= wdata[31:0];
end


//jump_type219
assign jump_type219_reg[31:0]   = jump_type219                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type219 <= 32'h0;
    else if( jump_type219_wr )
        jump_type219 <= wdata[31:0];
end


//jump_type220
assign jump_type220_reg[31:0]   = jump_type220                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type220 <= 32'h0;
    else if( jump_type220_wr )
        jump_type220 <= wdata[31:0];
end


//jump_type221
assign jump_type221_reg[31:0]   = jump_type221                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type221 <= 32'h0;
    else if( jump_type221_wr )
        jump_type221 <= wdata[31:0];
end


//jump_type222
assign jump_type222_reg[31:0]   = jump_type222                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type222 <= 32'h0;
    else if( jump_type222_wr )
        jump_type222 <= wdata[31:0];
end


//jump_type223
assign jump_type223_reg[31:0]   = jump_type223                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type223 <= 32'h0;
    else if( jump_type223_wr )
        jump_type223 <= wdata[31:0];
end


//jump_type224
assign jump_type224_reg[31:0]   = jump_type224                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type224 <= 32'h0;
    else if( jump_type224_wr )
        jump_type224 <= wdata[31:0];
end


//jump_type225
assign jump_type225_reg[31:0]   = jump_type225                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type225 <= 32'h0;
    else if( jump_type225_wr )
        jump_type225 <= wdata[31:0];
end


//jump_type226
assign jump_type226_reg[31:0]   = jump_type226                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type226 <= 32'h0;
    else if( jump_type226_wr )
        jump_type226 <= wdata[31:0];
end


//jump_type227
assign jump_type227_reg[31:0]   = jump_type227                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type227 <= 32'h0;
    else if( jump_type227_wr )
        jump_type227 <= wdata[31:0];
end


//jump_type228
assign jump_type228_reg[31:0]   = jump_type228                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type228 <= 32'h0;
    else if( jump_type228_wr )
        jump_type228 <= wdata[31:0];
end


//jump_type229
assign jump_type229_reg[31:0]   = jump_type229                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type229 <= 32'h0;
    else if( jump_type229_wr )
        jump_type229 <= wdata[31:0];
end


//jump_type230
assign jump_type230_reg[31:0]   = jump_type230                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type230 <= 32'h0;
    else if( jump_type230_wr )
        jump_type230 <= wdata[31:0];
end


//jump_type231
assign jump_type231_reg[31:0]   = jump_type231                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type231 <= 32'h0;
    else if( jump_type231_wr )
        jump_type231 <= wdata[31:0];
end


//jump_type232
assign jump_type232_reg[31:0]   = jump_type232                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type232 <= 32'h0;
    else if( jump_type232_wr )
        jump_type232 <= wdata[31:0];
end


//jump_type233
assign jump_type233_reg[31:0]   = jump_type233                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type233 <= 32'h0;
    else if( jump_type233_wr )
        jump_type233 <= wdata[31:0];
end


//jump_type234
assign jump_type234_reg[31:0]   = jump_type234                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type234 <= 32'h0;
    else if( jump_type234_wr )
        jump_type234 <= wdata[31:0];
end


//jump_type235
assign jump_type235_reg[31:0]   = jump_type235                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type235 <= 32'h0;
    else if( jump_type235_wr )
        jump_type235 <= wdata[31:0];
end


//jump_type236
assign jump_type236_reg[31:0]   = jump_type236                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type236 <= 32'h0;
    else if( jump_type236_wr )
        jump_type236 <= wdata[31:0];
end


//jump_type237
assign jump_type237_reg[31:0]   = jump_type237                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type237 <= 32'h0;
    else if( jump_type237_wr )
        jump_type237 <= wdata[31:0];
end


//jump_type238
assign jump_type238_reg[31:0]   = jump_type238                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type238 <= 32'h0;
    else if( jump_type238_wr )
        jump_type238 <= wdata[31:0];
end


//jump_type239
assign jump_type239_reg[31:0]   = jump_type239                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type239 <= 32'h0;
    else if( jump_type239_wr )
        jump_type239 <= wdata[31:0];
end


//jump_type240
assign jump_type240_reg[31:0]   = jump_type240                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type240 <= 32'h0;
    else if( jump_type240_wr )
        jump_type240 <= wdata[31:0];
end


//jump_type241
assign jump_type241_reg[31:0]   = jump_type241                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type241 <= 32'h0;
    else if( jump_type241_wr )
        jump_type241 <= wdata[31:0];
end


//jump_type242
assign jump_type242_reg[31:0]   = jump_type242                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type242 <= 32'h0;
    else if( jump_type242_wr )
        jump_type242 <= wdata[31:0];
end


//jump_type243
assign jump_type243_reg[31:0]   = jump_type243                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type243 <= 32'h0;
    else if( jump_type243_wr )
        jump_type243 <= wdata[31:0];
end


//jump_type244
assign jump_type244_reg[31:0]   = jump_type244                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type244 <= 32'h0;
    else if( jump_type244_wr )
        jump_type244 <= wdata[31:0];
end


//jump_type245
assign jump_type245_reg[31:0]   = jump_type245                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type245 <= 32'h0;
    else if( jump_type245_wr )
        jump_type245 <= wdata[31:0];
end


//jump_type246
assign jump_type246_reg[31:0]   = jump_type246                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type246 <= 32'h0;
    else if( jump_type246_wr )
        jump_type246 <= wdata[31:0];
end


//jump_type247
assign jump_type247_reg[31:0]   = jump_type247                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type247 <= 32'h0;
    else if( jump_type247_wr )
        jump_type247 <= wdata[31:0];
end


//jump_type248
assign jump_type248_reg[31:0]   = jump_type248                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type248 <= 32'h0;
    else if( jump_type248_wr )
        jump_type248 <= wdata[31:0];
end


//jump_type249
assign jump_type249_reg[31:0]   = jump_type249                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type249 <= 32'h0;
    else if( jump_type249_wr )
        jump_type249 <= wdata[31:0];
end


//jump_type250
assign jump_type250_reg[31:0]   = jump_type250                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type250 <= 32'h0;
    else if( jump_type250_wr )
        jump_type250 <= wdata[31:0];
end


//jump_type251
assign jump_type251_reg[31:0]   = jump_type251                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type251 <= 32'h0;
    else if( jump_type251_wr )
        jump_type251 <= wdata[31:0];
end


//jump_type252
assign jump_type252_reg[31:0]   = jump_type252                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type252 <= 32'h0;
    else if( jump_type252_wr )
        jump_type252 <= wdata[31:0];
end


//jump_type253
assign jump_type253_reg[31:0]   = jump_type253                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type253 <= 32'h0;
    else if( jump_type253_wr )
        jump_type253 <= wdata[31:0];
end


//jump_type254
assign jump_type254_reg[31:0]   = jump_type254                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type254 <= 32'h0;
    else if( jump_type254_wr )
        jump_type254 <= wdata[31:0];
end


//jump_type255
assign jump_type255_reg[31:0]   = jump_type255                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type255 <= 32'h0;
    else if( jump_type255_wr )
        jump_type255 <= wdata[31:0];
end


//jump_type256
assign jump_type256_reg[31:0]   = jump_type256                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type256 <= 32'h0;
    else if( jump_type256_wr )
        jump_type256 <= wdata[31:0];
end


//jump_type257
assign jump_type257_reg[31:0]   = jump_type257                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type257 <= 32'h0;
    else if( jump_type257_wr )
        jump_type257 <= wdata[31:0];
end


//jump_type258
assign jump_type258_reg[31:0]   = jump_type258                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type258 <= 32'h0;
    else if( jump_type258_wr )
        jump_type258 <= wdata[31:0];
end


//jump_type259
assign jump_type259_reg[31:0]   = jump_type259                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type259 <= 32'h0;
    else if( jump_type259_wr )
        jump_type259 <= wdata[31:0];
end


//jump_type260
assign jump_type260_reg[31:0]   = jump_type260                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type260 <= 32'h0;
    else if( jump_type260_wr )
        jump_type260 <= wdata[31:0];
end


//jump_type261
assign jump_type261_reg[31:0]   = jump_type261                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type261 <= 32'h0;
    else if( jump_type261_wr )
        jump_type261 <= wdata[31:0];
end


//jump_type262
assign jump_type262_reg[31:0]   = jump_type262                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type262 <= 32'h0;
    else if( jump_type262_wr )
        jump_type262 <= wdata[31:0];
end


//jump_type263
assign jump_type263_reg[31:0]   = jump_type263                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type263 <= 32'h0;
    else if( jump_type263_wr )
        jump_type263 <= wdata[31:0];
end


//jump_type264
assign jump_type264_reg[31:0]   = jump_type264                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type264 <= 32'h0;
    else if( jump_type264_wr )
        jump_type264 <= wdata[31:0];
end


//jump_type265
assign jump_type265_reg[31:0]   = jump_type265                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type265 <= 32'h0;
    else if( jump_type265_wr )
        jump_type265 <= wdata[31:0];
end


//jump_type266
assign jump_type266_reg[31:0]   = jump_type266                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type266 <= 32'h0;
    else if( jump_type266_wr )
        jump_type266 <= wdata[31:0];
end


//jump_type267
assign jump_type267_reg[31:0]   = jump_type267                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type267 <= 32'h0;
    else if( jump_type267_wr )
        jump_type267 <= wdata[31:0];
end


//jump_type268
assign jump_type268_reg[31:0]   = jump_type268                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type268 <= 32'h0;
    else if( jump_type268_wr )
        jump_type268 <= wdata[31:0];
end


//jump_type269
assign jump_type269_reg[31:0]   = jump_type269                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type269 <= 32'h0;
    else if( jump_type269_wr )
        jump_type269 <= wdata[31:0];
end


//jump_type270
assign jump_type270_reg[31:0]   = jump_type270                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type270 <= 32'h0;
    else if( jump_type270_wr )
        jump_type270 <= wdata[31:0];
end


//jump_type271
assign jump_type271_reg[31:0]   = jump_type271                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type271 <= 32'h0;
    else if( jump_type271_wr )
        jump_type271 <= wdata[31:0];
end


//jump_type272
assign jump_type272_reg[31:0]   = jump_type272                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type272 <= 32'h0;
    else if( jump_type272_wr )
        jump_type272 <= wdata[31:0];
end


//jump_type273
assign jump_type273_reg[31:0]   = jump_type273                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type273 <= 32'h0;
    else if( jump_type273_wr )
        jump_type273 <= wdata[31:0];
end


//jump_type274
assign jump_type274_reg[31:0]   = jump_type274                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type274 <= 32'h0;
    else if( jump_type274_wr )
        jump_type274 <= wdata[31:0];
end


//jump_type275
assign jump_type275_reg[31:0]   = jump_type275                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type275 <= 32'h0;
    else if( jump_type275_wr )
        jump_type275 <= wdata[31:0];
end


//jump_type276
assign jump_type276_reg[31:0]   = jump_type276                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type276 <= 32'h0;
    else if( jump_type276_wr )
        jump_type276 <= wdata[31:0];
end


//jump_type277
assign jump_type277_reg[31:0]   = jump_type277                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type277 <= 32'h0;
    else if( jump_type277_wr )
        jump_type277 <= wdata[31:0];
end


//jump_type278
assign jump_type278_reg[31:0]   = jump_type278                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type278 <= 32'h0;
    else if( jump_type278_wr )
        jump_type278 <= wdata[31:0];
end


//jump_type279
assign jump_type279_reg[31:0]   = jump_type279                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type279 <= 32'h0;
    else if( jump_type279_wr )
        jump_type279 <= wdata[31:0];
end


//jump_type280
assign jump_type280_reg[31:0]   = jump_type280                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type280 <= 32'h0;
    else if( jump_type280_wr )
        jump_type280 <= wdata[31:0];
end


//jump_type281
assign jump_type281_reg[31:0]   = jump_type281                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type281 <= 32'h0;
    else if( jump_type281_wr )
        jump_type281 <= wdata[31:0];
end


//jump_type282
assign jump_type282_reg[31:0]   = jump_type282                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type282 <= 32'h0;
    else if( jump_type282_wr )
        jump_type282 <= wdata[31:0];
end


//jump_type283
assign jump_type283_reg[31:0]   = jump_type283                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type283 <= 32'h0;
    else if( jump_type283_wr )
        jump_type283 <= wdata[31:0];
end


//jump_type284
assign jump_type284_reg[31:0]   = jump_type284                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type284 <= 32'h0;
    else if( jump_type284_wr )
        jump_type284 <= wdata[31:0];
end


//jump_type285
assign jump_type285_reg[31:0]   = jump_type285                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type285 <= 32'h0;
    else if( jump_type285_wr )
        jump_type285 <= wdata[31:0];
end


//jump_type286
assign jump_type286_reg[31:0]   = jump_type286                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type286 <= 32'h0;
    else if( jump_type286_wr )
        jump_type286 <= wdata[31:0];
end


//jump_type287
assign jump_type287_reg[31:0]   = jump_type287                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type287 <= 32'h0;
    else if( jump_type287_wr )
        jump_type287 <= wdata[31:0];
end


//jump_type288
assign jump_type288_reg[31:0]   = jump_type288                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type288 <= 32'h0;
    else if( jump_type288_wr )
        jump_type288 <= wdata[31:0];
end


//jump_type289
assign jump_type289_reg[31:0]   = jump_type289                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type289 <= 32'h0;
    else if( jump_type289_wr )
        jump_type289 <= wdata[31:0];
end


//jump_type290
assign jump_type290_reg[31:0]   = jump_type290                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type290 <= 32'h0;
    else if( jump_type290_wr )
        jump_type290 <= wdata[31:0];
end


//jump_type291
assign jump_type291_reg[31:0]   = jump_type291                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type291 <= 32'h0;
    else if( jump_type291_wr )
        jump_type291 <= wdata[31:0];
end


//jump_type292
assign jump_type292_reg[31:0]   = jump_type292                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type292 <= 32'h0;
    else if( jump_type292_wr )
        jump_type292 <= wdata[31:0];
end


//jump_type293
assign jump_type293_reg[31:0]   = jump_type293                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type293 <= 32'h0;
    else if( jump_type293_wr )
        jump_type293 <= wdata[31:0];
end


//jump_type294
assign jump_type294_reg[31:0]   = jump_type294                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type294 <= 32'h0;
    else if( jump_type294_wr )
        jump_type294 <= wdata[31:0];
end


//jump_type295
assign jump_type295_reg[31:0]   = jump_type295                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type295 <= 32'h0;
    else if( jump_type295_wr )
        jump_type295 <= wdata[31:0];
end


//jump_type296
assign jump_type296_reg[31:0]   = jump_type296                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type296 <= 32'h0;
    else if( jump_type296_wr )
        jump_type296 <= wdata[31:0];
end


//jump_type297
assign jump_type297_reg[31:0]   = jump_type297                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type297 <= 32'h0;
    else if( jump_type297_wr )
        jump_type297 <= wdata[31:0];
end


//jump_type298
assign jump_type298_reg[31:0]   = jump_type298                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type298 <= 32'h0;
    else if( jump_type298_wr )
        jump_type298 <= wdata[31:0];
end


//jump_type299
assign jump_type299_reg[31:0]   = jump_type299                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type299 <= 32'h0;
    else if( jump_type299_wr )
        jump_type299 <= wdata[31:0];
end


//jump_type300
assign jump_type300_reg[31:0]   = jump_type300                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type300 <= 32'h0;
    else if( jump_type300_wr )
        jump_type300 <= wdata[31:0];
end


//jump_type301
assign jump_type301_reg[31:0]   = jump_type301                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type301 <= 32'h0;
    else if( jump_type301_wr )
        jump_type301 <= wdata[31:0];
end


//jump_type302
assign jump_type302_reg[31:0]   = jump_type302                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type302 <= 32'h0;
    else if( jump_type302_wr )
        jump_type302 <= wdata[31:0];
end


//jump_type303
assign jump_type303_reg[31:0]   = jump_type303                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type303 <= 32'h0;
    else if( jump_type303_wr )
        jump_type303 <= wdata[31:0];
end


//jump_type304
assign jump_type304_reg[31:0]   = jump_type304                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type304 <= 32'h0;
    else if( jump_type304_wr )
        jump_type304 <= wdata[31:0];
end


//jump_type305
assign jump_type305_reg[31:0]   = jump_type305                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type305 <= 32'h0;
    else if( jump_type305_wr )
        jump_type305 <= wdata[31:0];
end


//jump_type306
assign jump_type306_reg[31:0]   = jump_type306                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type306 <= 32'h0;
    else if( jump_type306_wr )
        jump_type306 <= wdata[31:0];
end


//jump_type307
assign jump_type307_reg[31:0]   = jump_type307                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type307 <= 32'h0;
    else if( jump_type307_wr )
        jump_type307 <= wdata[31:0];
end


//jump_type308
assign jump_type308_reg[31:0]   = jump_type308                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type308 <= 32'h0;
    else if( jump_type308_wr )
        jump_type308 <= wdata[31:0];
end


//jump_type309
assign jump_type309_reg[31:0]   = jump_type309                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type309 <= 32'h0;
    else if( jump_type309_wr )
        jump_type309 <= wdata[31:0];
end


//jump_type310
assign jump_type310_reg[31:0]   = jump_type310                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type310 <= 32'h0;
    else if( jump_type310_wr )
        jump_type310 <= wdata[31:0];
end


//jump_type311
assign jump_type311_reg[31:0]   = jump_type311                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type311 <= 32'h0;
    else if( jump_type311_wr )
        jump_type311 <= wdata[31:0];
end


//jump_type312
assign jump_type312_reg[31:0]   = jump_type312                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type312 <= 32'h0;
    else if( jump_type312_wr )
        jump_type312 <= wdata[31:0];
end


//jump_type313
assign jump_type313_reg[31:0]   = jump_type313                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type313 <= 32'h0;
    else if( jump_type313_wr )
        jump_type313 <= wdata[31:0];
end


//jump_type314
assign jump_type314_reg[31:0]   = jump_type314                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type314 <= 32'h0;
    else if( jump_type314_wr )
        jump_type314 <= wdata[31:0];
end


//jump_type315
assign jump_type315_reg[31:0]   = jump_type315                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type315 <= 32'h0;
    else if( jump_type315_wr )
        jump_type315 <= wdata[31:0];
end


//jump_type316
assign jump_type316_reg[31:0]   = jump_type316                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type316 <= 32'h0;
    else if( jump_type316_wr )
        jump_type316 <= wdata[31:0];
end


//jump_type317
assign jump_type317_reg[31:0]   = jump_type317                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type317 <= 32'h0;
    else if( jump_type317_wr )
        jump_type317 <= wdata[31:0];
end


//jump_type318
assign jump_type318_reg[31:0]   = jump_type318                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type318 <= 32'h0;
    else if( jump_type318_wr )
        jump_type318 <= wdata[31:0];
end


//jump_type319
assign jump_type319_reg[31:0]   = jump_type319                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type319 <= 32'h0;
    else if( jump_type319_wr )
        jump_type319 <= wdata[31:0];
end


//jump_type320
assign jump_type320_reg[31:0]   = jump_type320                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type320 <= 32'h0;
    else if( jump_type320_wr )
        jump_type320 <= wdata[31:0];
end


//jump_type321
assign jump_type321_reg[31:0]   = jump_type321                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type321 <= 32'h0;
    else if( jump_type321_wr )
        jump_type321 <= wdata[31:0];
end


//jump_type322
assign jump_type322_reg[31:0]   = jump_type322                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type322 <= 32'h0;
    else if( jump_type322_wr )
        jump_type322 <= wdata[31:0];
end


//jump_type323
assign jump_type323_reg[31:0]   = jump_type323                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type323 <= 32'h0;
    else if( jump_type323_wr )
        jump_type323 <= wdata[31:0];
end


//jump_type324
assign jump_type324_reg[31:0]   = jump_type324                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type324 <= 32'h0;
    else if( jump_type324_wr )
        jump_type324 <= wdata[31:0];
end


//jump_type325
assign jump_type325_reg[31:0]   = jump_type325                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type325 <= 32'h0;
    else if( jump_type325_wr )
        jump_type325 <= wdata[31:0];
end


//jump_type326
assign jump_type326_reg[31:0]   = jump_type326                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type326 <= 32'h0;
    else if( jump_type326_wr )
        jump_type326 <= wdata[31:0];
end


//jump_type327
assign jump_type327_reg[31:0]   = jump_type327                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type327 <= 32'h0;
    else if( jump_type327_wr )
        jump_type327 <= wdata[31:0];
end


//jump_type328
assign jump_type328_reg[31:0]   = jump_type328                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type328 <= 32'h0;
    else if( jump_type328_wr )
        jump_type328 <= wdata[31:0];
end


//jump_type329
assign jump_type329_reg[31:0]   = jump_type329                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type329 <= 32'h0;
    else if( jump_type329_wr )
        jump_type329 <= wdata[31:0];
end


//jump_type330
assign jump_type330_reg[31:0]   = jump_type330                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type330 <= 32'h0;
    else if( jump_type330_wr )
        jump_type330 <= wdata[31:0];
end


//jump_type331
assign jump_type331_reg[31:0]   = jump_type331                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type331 <= 32'h0;
    else if( jump_type331_wr )
        jump_type331 <= wdata[31:0];
end


//jump_type332
assign jump_type332_reg[31:0]   = jump_type332                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type332 <= 32'h0;
    else if( jump_type332_wr )
        jump_type332 <= wdata[31:0];
end


//jump_type333
assign jump_type333_reg[31:0]   = jump_type333                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type333 <= 32'h0;
    else if( jump_type333_wr )
        jump_type333 <= wdata[31:0];
end


//jump_type334
assign jump_type334_reg[31:0]   = jump_type334                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type334 <= 32'h0;
    else if( jump_type334_wr )
        jump_type334 <= wdata[31:0];
end


//jump_type335
assign jump_type335_reg[31:0]   = jump_type335                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type335 <= 32'h0;
    else if( jump_type335_wr )
        jump_type335 <= wdata[31:0];
end


//jump_type336
assign jump_type336_reg[31:0]   = jump_type336                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type336 <= 32'h0;
    else if( jump_type336_wr )
        jump_type336 <= wdata[31:0];
end


//jump_type337
assign jump_type337_reg[31:0]   = jump_type337                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type337 <= 32'h0;
    else if( jump_type337_wr )
        jump_type337 <= wdata[31:0];
end


//jump_type338
assign jump_type338_reg[31:0]   = jump_type338                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type338 <= 32'h0;
    else if( jump_type338_wr )
        jump_type338 <= wdata[31:0];
end


//jump_type339
assign jump_type339_reg[31:0]   = jump_type339                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type339 <= 32'h0;
    else if( jump_type339_wr )
        jump_type339 <= wdata[31:0];
end


//jump_type340
assign jump_type340_reg[31:0]   = jump_type340                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type340 <= 32'h0;
    else if( jump_type340_wr )
        jump_type340 <= wdata[31:0];
end


//jump_type341
assign jump_type341_reg[31:0]   = jump_type341                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type341 <= 32'h0;
    else if( jump_type341_wr )
        jump_type341 <= wdata[31:0];
end


//jump_type342
assign jump_type342_reg[31:0]   = jump_type342                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type342 <= 32'h0;
    else if( jump_type342_wr )
        jump_type342 <= wdata[31:0];
end


//jump_type343
assign jump_type343_reg[31:0]   = jump_type343                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type343 <= 32'h0;
    else if( jump_type343_wr )
        jump_type343 <= wdata[31:0];
end


//jump_type344
assign jump_type344_reg[31:0]   = jump_type344                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type344 <= 32'h0;
    else if( jump_type344_wr )
        jump_type344 <= wdata[31:0];
end


//jump_type345
assign jump_type345_reg[31:0]   = jump_type345                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type345 <= 32'h0;
    else if( jump_type345_wr )
        jump_type345 <= wdata[31:0];
end


//jump_type346
assign jump_type346_reg[31:0]   = jump_type346                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type346 <= 32'h0;
    else if( jump_type346_wr )
        jump_type346 <= wdata[31:0];
end


//jump_type347
assign jump_type347_reg[31:0]   = jump_type347                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type347 <= 32'h0;
    else if( jump_type347_wr )
        jump_type347 <= wdata[31:0];
end


//jump_type348
assign jump_type348_reg[31:0]   = jump_type348                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type348 <= 32'h0;
    else if( jump_type348_wr )
        jump_type348 <= wdata[31:0];
end


//jump_type349
assign jump_type349_reg[31:0]   = jump_type349                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type349 <= 32'h0;
    else if( jump_type349_wr )
        jump_type349 <= wdata[31:0];
end


//jump_type350
assign jump_type350_reg[31:0]   = jump_type350                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type350 <= 32'h0;
    else if( jump_type350_wr )
        jump_type350 <= wdata[31:0];
end


//jump_type351
assign jump_type351_reg[31:0]   = jump_type351                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type351 <= 32'h0;
    else if( jump_type351_wr )
        jump_type351 <= wdata[31:0];
end


//jump_type352
assign jump_type352_reg[31:0]   = jump_type352                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type352 <= 32'h0;
    else if( jump_type352_wr )
        jump_type352 <= wdata[31:0];
end


//jump_type353
assign jump_type353_reg[31:0]   = jump_type353                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type353 <= 32'h0;
    else if( jump_type353_wr )
        jump_type353 <= wdata[31:0];
end


//jump_type354
assign jump_type354_reg[31:0]   = jump_type354                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type354 <= 32'h0;
    else if( jump_type354_wr )
        jump_type354 <= wdata[31:0];
end


//jump_type355
assign jump_type355_reg[31:0]   = jump_type355                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type355 <= 32'h0;
    else if( jump_type355_wr )
        jump_type355 <= wdata[31:0];
end


//jump_type356
assign jump_type356_reg[31:0]   = jump_type356                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type356 <= 32'h0;
    else if( jump_type356_wr )
        jump_type356 <= wdata[31:0];
end


//jump_type357
assign jump_type357_reg[31:0]   = jump_type357                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type357 <= 32'h0;
    else if( jump_type357_wr )
        jump_type357 <= wdata[31:0];
end


//jump_type358
assign jump_type358_reg[31:0]   = jump_type358                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type358 <= 32'h0;
    else if( jump_type358_wr )
        jump_type358 <= wdata[31:0];
end


//jump_type359
assign jump_type359_reg[31:0]   = jump_type359                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type359 <= 32'h0;
    else if( jump_type359_wr )
        jump_type359 <= wdata[31:0];
end


//jump_type360
assign jump_type360_reg[31:0]   = jump_type360                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type360 <= 32'h0;
    else if( jump_type360_wr )
        jump_type360 <= wdata[31:0];
end


//jump_type361
assign jump_type361_reg[31:0]   = jump_type361                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type361 <= 32'h0;
    else if( jump_type361_wr )
        jump_type361 <= wdata[31:0];
end


//jump_type362
assign jump_type362_reg[31:0]   = jump_type362                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type362 <= 32'h0;
    else if( jump_type362_wr )
        jump_type362 <= wdata[31:0];
end


//jump_type363
assign jump_type363_reg[31:0]   = jump_type363                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type363 <= 32'h0;
    else if( jump_type363_wr )
        jump_type363 <= wdata[31:0];
end


//jump_type364
assign jump_type364_reg[31:0]   = jump_type364                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type364 <= 32'h0;
    else if( jump_type364_wr )
        jump_type364 <= wdata[31:0];
end


//jump_type365
assign jump_type365_reg[31:0]   = jump_type365                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type365 <= 32'h0;
    else if( jump_type365_wr )
        jump_type365 <= wdata[31:0];
end


//jump_type366
assign jump_type366_reg[31:0]   = jump_type366                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type366 <= 32'h0;
    else if( jump_type366_wr )
        jump_type366 <= wdata[31:0];
end


//jump_type367
assign jump_type367_reg[31:0]   = jump_type367                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type367 <= 32'h0;
    else if( jump_type367_wr )
        jump_type367 <= wdata[31:0];
end


//jump_type368
assign jump_type368_reg[31:0]   = jump_type368                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type368 <= 32'h0;
    else if( jump_type368_wr )
        jump_type368 <= wdata[31:0];
end


//jump_type369
assign jump_type369_reg[31:0]   = jump_type369                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type369 <= 32'h0;
    else if( jump_type369_wr )
        jump_type369 <= wdata[31:0];
end


//jump_type370
assign jump_type370_reg[31:0]   = jump_type370                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type370 <= 32'h0;
    else if( jump_type370_wr )
        jump_type370 <= wdata[31:0];
end


//jump_type371
assign jump_type371_reg[31:0]   = jump_type371                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type371 <= 32'h0;
    else if( jump_type371_wr )
        jump_type371 <= wdata[31:0];
end


//jump_type372
assign jump_type372_reg[31:0]   = jump_type372                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type372 <= 32'h0;
    else if( jump_type372_wr )
        jump_type372 <= wdata[31:0];
end


//jump_type373
assign jump_type373_reg[31:0]   = jump_type373                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type373 <= 32'h0;
    else if( jump_type373_wr )
        jump_type373 <= wdata[31:0];
end


//jump_type374
assign jump_type374_reg[31:0]   = jump_type374                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type374 <= 32'h0;
    else if( jump_type374_wr )
        jump_type374 <= wdata[31:0];
end


//jump_type375
assign jump_type375_reg[31:0]   = jump_type375                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type375 <= 32'h0;
    else if( jump_type375_wr )
        jump_type375 <= wdata[31:0];
end


//jump_type376
assign jump_type376_reg[31:0]   = jump_type376                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type376 <= 32'h0;
    else if( jump_type376_wr )
        jump_type376 <= wdata[31:0];
end


//jump_type377
assign jump_type377_reg[31:0]   = jump_type377                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type377 <= 32'h0;
    else if( jump_type377_wr )
        jump_type377 <= wdata[31:0];
end


//jump_type378
assign jump_type378_reg[31:0]   = jump_type378                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type378 <= 32'h0;
    else if( jump_type378_wr )
        jump_type378 <= wdata[31:0];
end


//jump_type379
assign jump_type379_reg[31:0]   = jump_type379                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type379 <= 32'h0;
    else if( jump_type379_wr )
        jump_type379 <= wdata[31:0];
end


//jump_type380
assign jump_type380_reg[31:0]   = jump_type380                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type380 <= 32'h0;
    else if( jump_type380_wr )
        jump_type380 <= wdata[31:0];
end


//jump_type381
assign jump_type381_reg[31:0]   = jump_type381                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type381 <= 32'h0;
    else if( jump_type381_wr )
        jump_type381 <= wdata[31:0];
end


//jump_type382
assign jump_type382_reg[31:0]   = jump_type382                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type382 <= 32'h0;
    else if( jump_type382_wr )
        jump_type382 <= wdata[31:0];
end


//jump_type383
assign jump_type383_reg[31:0]   = jump_type383                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type383 <= 32'h0;
    else if( jump_type383_wr )
        jump_type383 <= wdata[31:0];
end


//jump_type384
assign jump_type384_reg[31:0]   = jump_type384                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type384 <= 32'h0;
    else if( jump_type384_wr )
        jump_type384 <= wdata[31:0];
end


//jump_type385
assign jump_type385_reg[31:0]   = jump_type385                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type385 <= 32'h0;
    else if( jump_type385_wr )
        jump_type385 <= wdata[31:0];
end


//jump_type386
assign jump_type386_reg[31:0]   = jump_type386                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type386 <= 32'h0;
    else if( jump_type386_wr )
        jump_type386 <= wdata[31:0];
end


//jump_type387
assign jump_type387_reg[31:0]   = jump_type387                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type387 <= 32'h0;
    else if( jump_type387_wr )
        jump_type387 <= wdata[31:0];
end


//jump_type388
assign jump_type388_reg[31:0]   = jump_type388                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type388 <= 32'h0;
    else if( jump_type388_wr )
        jump_type388 <= wdata[31:0];
end


//jump_type389
assign jump_type389_reg[31:0]   = jump_type389                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type389 <= 32'h0;
    else if( jump_type389_wr )
        jump_type389 <= wdata[31:0];
end


//jump_type390
assign jump_type390_reg[31:0]   = jump_type390                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type390 <= 32'h0;
    else if( jump_type390_wr )
        jump_type390 <= wdata[31:0];
end


//jump_type391
assign jump_type391_reg[31:0]   = jump_type391                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type391 <= 32'h0;
    else if( jump_type391_wr )
        jump_type391 <= wdata[31:0];
end


//jump_type392
assign jump_type392_reg[31:0]   = jump_type392                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type392 <= 32'h0;
    else if( jump_type392_wr )
        jump_type392 <= wdata[31:0];
end


//jump_type393
assign jump_type393_reg[31:0]   = jump_type393                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type393 <= 32'h0;
    else if( jump_type393_wr )
        jump_type393 <= wdata[31:0];
end


//jump_type394
assign jump_type394_reg[31:0]   = jump_type394                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type394 <= 32'h0;
    else if( jump_type394_wr )
        jump_type394 <= wdata[31:0];
end


//jump_type395
assign jump_type395_reg[31:0]   = jump_type395                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type395 <= 32'h0;
    else if( jump_type395_wr )
        jump_type395 <= wdata[31:0];
end


//jump_type396
assign jump_type396_reg[31:0]   = jump_type396                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type396 <= 32'h0;
    else if( jump_type396_wr )
        jump_type396 <= wdata[31:0];
end


//jump_type397
assign jump_type397_reg[31:0]   = jump_type397                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type397 <= 32'h0;
    else if( jump_type397_wr )
        jump_type397 <= wdata[31:0];
end


//jump_type398
assign jump_type398_reg[31:0]   = jump_type398                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type398 <= 32'h0;
    else if( jump_type398_wr )
        jump_type398 <= wdata[31:0];
end


//jump_type399
assign jump_type399_reg[31:0]   = jump_type399                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type399 <= 32'h0;
    else if( jump_type399_wr )
        jump_type399 <= wdata[31:0];
end


//jump_type400
assign jump_type400_reg[31:0]   = jump_type400                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type400 <= 32'h0;
    else if( jump_type400_wr )
        jump_type400 <= wdata[31:0];
end


//jump_type401
assign jump_type401_reg[31:0]   = jump_type401                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type401 <= 32'h0;
    else if( jump_type401_wr )
        jump_type401 <= wdata[31:0];
end


//jump_type402
assign jump_type402_reg[31:0]   = jump_type402                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type402 <= 32'h0;
    else if( jump_type402_wr )
        jump_type402 <= wdata[31:0];
end


//jump_type403
assign jump_type403_reg[31:0]   = jump_type403                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type403 <= 32'h0;
    else if( jump_type403_wr )
        jump_type403 <= wdata[31:0];
end


//jump_type404
assign jump_type404_reg[31:0]   = jump_type404                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type404 <= 32'h0;
    else if( jump_type404_wr )
        jump_type404 <= wdata[31:0];
end


//jump_type405
assign jump_type405_reg[31:0]   = jump_type405                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type405 <= 32'h0;
    else if( jump_type405_wr )
        jump_type405 <= wdata[31:0];
end


//jump_type406
assign jump_type406_reg[31:0]   = jump_type406                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type406 <= 32'h0;
    else if( jump_type406_wr )
        jump_type406 <= wdata[31:0];
end


//jump_type407
assign jump_type407_reg[31:0]   = jump_type407                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type407 <= 32'h0;
    else if( jump_type407_wr )
        jump_type407 <= wdata[31:0];
end


//jump_type408
assign jump_type408_reg[31:0]   = jump_type408                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type408 <= 32'h0;
    else if( jump_type408_wr )
        jump_type408 <= wdata[31:0];
end


//jump_type409
assign jump_type409_reg[31:0]   = jump_type409                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type409 <= 32'h0;
    else if( jump_type409_wr )
        jump_type409 <= wdata[31:0];
end


//jump_type410
assign jump_type410_reg[31:0]   = jump_type410                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type410 <= 32'h0;
    else if( jump_type410_wr )
        jump_type410 <= wdata[31:0];
end


//jump_type411
assign jump_type411_reg[31:0]   = jump_type411                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type411 <= 32'h0;
    else if( jump_type411_wr )
        jump_type411 <= wdata[31:0];
end


//jump_type412
assign jump_type412_reg[31:0]   = jump_type412                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type412 <= 32'h0;
    else if( jump_type412_wr )
        jump_type412 <= wdata[31:0];
end


//jump_type413
assign jump_type413_reg[31:0]   = jump_type413                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type413 <= 32'h0;
    else if( jump_type413_wr )
        jump_type413 <= wdata[31:0];
end


//jump_type414
assign jump_type414_reg[31:0]   = jump_type414                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type414 <= 32'h0;
    else if( jump_type414_wr )
        jump_type414 <= wdata[31:0];
end


//jump_type415
assign jump_type415_reg[31:0]   = jump_type415                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type415 <= 32'h0;
    else if( jump_type415_wr )
        jump_type415 <= wdata[31:0];
end


//jump_type416
assign jump_type416_reg[31:0]   = jump_type416                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type416 <= 32'h0;
    else if( jump_type416_wr )
        jump_type416 <= wdata[31:0];
end


//jump_type417
assign jump_type417_reg[31:0]   = jump_type417                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type417 <= 32'h0;
    else if( jump_type417_wr )
        jump_type417 <= wdata[31:0];
end


//jump_type418
assign jump_type418_reg[31:0]   = jump_type418                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type418 <= 32'h0;
    else if( jump_type418_wr )
        jump_type418 <= wdata[31:0];
end


//jump_type419
assign jump_type419_reg[31:0]   = jump_type419                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type419 <= 32'h0;
    else if( jump_type419_wr )
        jump_type419 <= wdata[31:0];
end


//jump_type420
assign jump_type420_reg[31:0]   = jump_type420                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type420 <= 32'h0;
    else if( jump_type420_wr )
        jump_type420 <= wdata[31:0];
end


//jump_type421
assign jump_type421_reg[31:0]   = jump_type421                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type421 <= 32'h0;
    else if( jump_type421_wr )
        jump_type421 <= wdata[31:0];
end


//jump_type422
assign jump_type422_reg[31:0]   = jump_type422                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type422 <= 32'h0;
    else if( jump_type422_wr )
        jump_type422 <= wdata[31:0];
end


//jump_type423
assign jump_type423_reg[31:0]   = jump_type423                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type423 <= 32'h0;
    else if( jump_type423_wr )
        jump_type423 <= wdata[31:0];
end


//jump_type424
assign jump_type424_reg[31:0]   = jump_type424                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type424 <= 32'h0;
    else if( jump_type424_wr )
        jump_type424 <= wdata[31:0];
end


//jump_type425
assign jump_type425_reg[31:0]   = jump_type425                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type425 <= 32'h0;
    else if( jump_type425_wr )
        jump_type425 <= wdata[31:0];
end


//jump_type426
assign jump_type426_reg[31:0]   = jump_type426                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type426 <= 32'h0;
    else if( jump_type426_wr )
        jump_type426 <= wdata[31:0];
end


//jump_type427
assign jump_type427_reg[31:0]   = jump_type427                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type427 <= 32'h0;
    else if( jump_type427_wr )
        jump_type427 <= wdata[31:0];
end


//jump_type428
assign jump_type428_reg[31:0]   = jump_type428                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type428 <= 32'h0;
    else if( jump_type428_wr )
        jump_type428 <= wdata[31:0];
end


//jump_type429
assign jump_type429_reg[31:0]   = jump_type429                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type429 <= 32'h0;
    else if( jump_type429_wr )
        jump_type429 <= wdata[31:0];
end


//jump_type430
assign jump_type430_reg[31:0]   = jump_type430                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type430 <= 32'h0;
    else if( jump_type430_wr )
        jump_type430 <= wdata[31:0];
end


//jump_type431
assign jump_type431_reg[31:0]   = jump_type431                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type431 <= 32'h0;
    else if( jump_type431_wr )
        jump_type431 <= wdata[31:0];
end


//jump_type432
assign jump_type432_reg[31:0]   = jump_type432                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type432 <= 32'h0;
    else if( jump_type432_wr )
        jump_type432 <= wdata[31:0];
end


//jump_type433
assign jump_type433_reg[31:0]   = jump_type433                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type433 <= 32'h0;
    else if( jump_type433_wr )
        jump_type433 <= wdata[31:0];
end


//jump_type434
assign jump_type434_reg[31:0]   = jump_type434                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type434 <= 32'h0;
    else if( jump_type434_wr )
        jump_type434 <= wdata[31:0];
end


//jump_type435
assign jump_type435_reg[31:0]   = jump_type435                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type435 <= 32'h0;
    else if( jump_type435_wr )
        jump_type435 <= wdata[31:0];
end


//jump_type436
assign jump_type436_reg[31:0]   = jump_type436                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type436 <= 32'h0;
    else if( jump_type436_wr )
        jump_type436 <= wdata[31:0];
end


//jump_type437
assign jump_type437_reg[31:0]   = jump_type437                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type437 <= 32'h0;
    else if( jump_type437_wr )
        jump_type437 <= wdata[31:0];
end


//jump_type438
assign jump_type438_reg[31:0]   = jump_type438                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type438 <= 32'h0;
    else if( jump_type438_wr )
        jump_type438 <= wdata[31:0];
end


//jump_type439
assign jump_type439_reg[31:0]   = jump_type439                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type439 <= 32'h0;
    else if( jump_type439_wr )
        jump_type439 <= wdata[31:0];
end


//jump_type440
assign jump_type440_reg[31:0]   = jump_type440                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type440 <= 32'h0;
    else if( jump_type440_wr )
        jump_type440 <= wdata[31:0];
end


//jump_type441
assign jump_type441_reg[31:0]   = jump_type441                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type441 <= 32'h0;
    else if( jump_type441_wr )
        jump_type441 <= wdata[31:0];
end


//jump_type442
assign jump_type442_reg[31:0]   = jump_type442                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type442 <= 32'h0;
    else if( jump_type442_wr )
        jump_type442 <= wdata[31:0];
end


//jump_type443
assign jump_type443_reg[31:0]   = jump_type443                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type443 <= 32'h0;
    else if( jump_type443_wr )
        jump_type443 <= wdata[31:0];
end


//jump_type444
assign jump_type444_reg[31:0]   = jump_type444                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type444 <= 32'h0;
    else if( jump_type444_wr )
        jump_type444 <= wdata[31:0];
end


//jump_type445
assign jump_type445_reg[31:0]   = jump_type445                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type445 <= 32'h0;
    else if( jump_type445_wr )
        jump_type445 <= wdata[31:0];
end


//jump_type446
assign jump_type446_reg[31:0]   = jump_type446                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type446 <= 32'h0;
    else if( jump_type446_wr )
        jump_type446 <= wdata[31:0];
end


//jump_type447
assign jump_type447_reg[31:0]   = jump_type447                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type447 <= 32'h0;
    else if( jump_type447_wr )
        jump_type447 <= wdata[31:0];
end


//jump_type448
assign jump_type448_reg[31:0]   = jump_type448                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type448 <= 32'h0;
    else if( jump_type448_wr )
        jump_type448 <= wdata[31:0];
end


//jump_type449
assign jump_type449_reg[31:0]   = jump_type449                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type449 <= 32'h0;
    else if( jump_type449_wr )
        jump_type449 <= wdata[31:0];
end


//jump_type450
assign jump_type450_reg[31:0]   = jump_type450                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type450 <= 32'h0;
    else if( jump_type450_wr )
        jump_type450 <= wdata[31:0];
end


//jump_type451
assign jump_type451_reg[31:0]   = jump_type451                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type451 <= 32'h0;
    else if( jump_type451_wr )
        jump_type451 <= wdata[31:0];
end


//jump_type452
assign jump_type452_reg[31:0]   = jump_type452                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type452 <= 32'h0;
    else if( jump_type452_wr )
        jump_type452 <= wdata[31:0];
end


//jump_type453
assign jump_type453_reg[31:0]   = jump_type453                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type453 <= 32'h0;
    else if( jump_type453_wr )
        jump_type453 <= wdata[31:0];
end


//jump_type454
assign jump_type454_reg[31:0]   = jump_type454                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type454 <= 32'h0;
    else if( jump_type454_wr )
        jump_type454 <= wdata[31:0];
end


//jump_type455
assign jump_type455_reg[31:0]   = jump_type455                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type455 <= 32'h0;
    else if( jump_type455_wr )
        jump_type455 <= wdata[31:0];
end


//jump_type456
assign jump_type456_reg[31:0]   = jump_type456                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type456 <= 32'h0;
    else if( jump_type456_wr )
        jump_type456 <= wdata[31:0];
end


//jump_type457
assign jump_type457_reg[31:0]   = jump_type457                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type457 <= 32'h0;
    else if( jump_type457_wr )
        jump_type457 <= wdata[31:0];
end


//jump_type458
assign jump_type458_reg[31:0]   = jump_type458                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type458 <= 32'h0;
    else if( jump_type458_wr )
        jump_type458 <= wdata[31:0];
end


//jump_type459
assign jump_type459_reg[31:0]   = jump_type459                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type459 <= 32'h0;
    else if( jump_type459_wr )
        jump_type459 <= wdata[31:0];
end


//jump_type460
assign jump_type460_reg[31:0]   = jump_type460                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type460 <= 32'h0;
    else if( jump_type460_wr )
        jump_type460 <= wdata[31:0];
end


//jump_type461
assign jump_type461_reg[31:0]   = jump_type461                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type461 <= 32'h0;
    else if( jump_type461_wr )
        jump_type461 <= wdata[31:0];
end


//jump_type462
assign jump_type462_reg[31:0]   = jump_type462                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type462 <= 32'h0;
    else if( jump_type462_wr )
        jump_type462 <= wdata[31:0];
end


//jump_type463
assign jump_type463_reg[31:0]   = jump_type463                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type463 <= 32'h0;
    else if( jump_type463_wr )
        jump_type463 <= wdata[31:0];
end


//jump_type464
assign jump_type464_reg[31:0]   = jump_type464                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type464 <= 32'h0;
    else if( jump_type464_wr )
        jump_type464 <= wdata[31:0];
end


//jump_type465
assign jump_type465_reg[31:0]   = jump_type465                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type465 <= 32'h0;
    else if( jump_type465_wr )
        jump_type465 <= wdata[31:0];
end


//jump_type466
assign jump_type466_reg[31:0]   = jump_type466                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type466 <= 32'h0;
    else if( jump_type466_wr )
        jump_type466 <= wdata[31:0];
end


//jump_type467
assign jump_type467_reg[31:0]   = jump_type467                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type467 <= 32'h0;
    else if( jump_type467_wr )
        jump_type467 <= wdata[31:0];
end


//jump_type468
assign jump_type468_reg[31:0]   = jump_type468                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type468 <= 32'h0;
    else if( jump_type468_wr )
        jump_type468 <= wdata[31:0];
end


//jump_type469
assign jump_type469_reg[31:0]   = jump_type469                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type469 <= 32'h0;
    else if( jump_type469_wr )
        jump_type469 <= wdata[31:0];
end


//jump_type470
assign jump_type470_reg[31:0]   = jump_type470                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type470 <= 32'h0;
    else if( jump_type470_wr )
        jump_type470 <= wdata[31:0];
end


//jump_type471
assign jump_type471_reg[31:0]   = jump_type471                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type471 <= 32'h0;
    else if( jump_type471_wr )
        jump_type471 <= wdata[31:0];
end


//jump_type472
assign jump_type472_reg[31:0]   = jump_type472                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type472 <= 32'h0;
    else if( jump_type472_wr )
        jump_type472 <= wdata[31:0];
end


//jump_type473
assign jump_type473_reg[31:0]   = jump_type473                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type473 <= 32'h0;
    else if( jump_type473_wr )
        jump_type473 <= wdata[31:0];
end


//jump_type474
assign jump_type474_reg[31:0]   = jump_type474                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type474 <= 32'h0;
    else if( jump_type474_wr )
        jump_type474 <= wdata[31:0];
end


//jump_type475
assign jump_type475_reg[31:0]   = jump_type475                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type475 <= 32'h0;
    else if( jump_type475_wr )
        jump_type475 <= wdata[31:0];
end


//jump_type476
assign jump_type476_reg[31:0]   = jump_type476                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type476 <= 32'h0;
    else if( jump_type476_wr )
        jump_type476 <= wdata[31:0];
end


//jump_type477
assign jump_type477_reg[31:0]   = jump_type477                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type477 <= 32'h0;
    else if( jump_type477_wr )
        jump_type477 <= wdata[31:0];
end


//jump_type478
assign jump_type478_reg[31:0]   = jump_type478                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type478 <= 32'h0;
    else if( jump_type478_wr )
        jump_type478 <= wdata[31:0];
end


//jump_type479
assign jump_type479_reg[31:0]   = jump_type479                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type479 <= 32'h0;
    else if( jump_type479_wr )
        jump_type479 <= wdata[31:0];
end


//jump_type480
assign jump_type480_reg[31:0]   = jump_type480                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type480 <= 32'h0;
    else if( jump_type480_wr )
        jump_type480 <= wdata[31:0];
end


//jump_type481
assign jump_type481_reg[31:0]   = jump_type481                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type481 <= 32'h0;
    else if( jump_type481_wr )
        jump_type481 <= wdata[31:0];
end


//jump_type482
assign jump_type482_reg[31:0]   = jump_type482                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type482 <= 32'h0;
    else if( jump_type482_wr )
        jump_type482 <= wdata[31:0];
end


//jump_type483
assign jump_type483_reg[31:0]   = jump_type483                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type483 <= 32'h0;
    else if( jump_type483_wr )
        jump_type483 <= wdata[31:0];
end


//jump_type484
assign jump_type484_reg[31:0]   = jump_type484                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type484 <= 32'h0;
    else if( jump_type484_wr )
        jump_type484 <= wdata[31:0];
end


//jump_type485
assign jump_type485_reg[31:0]   = jump_type485                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type485 <= 32'h0;
    else if( jump_type485_wr )
        jump_type485 <= wdata[31:0];
end


//jump_type486
assign jump_type486_reg[31:0]   = jump_type486                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type486 <= 32'h0;
    else if( jump_type486_wr )
        jump_type486 <= wdata[31:0];
end


//jump_type487
assign jump_type487_reg[31:0]   = jump_type487                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type487 <= 32'h0;
    else if( jump_type487_wr )
        jump_type487 <= wdata[31:0];
end


//jump_type488
assign jump_type488_reg[31:0]   = jump_type488                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type488 <= 32'h0;
    else if( jump_type488_wr )
        jump_type488 <= wdata[31:0];
end


//jump_type489
assign jump_type489_reg[31:0]   = jump_type489                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type489 <= 32'h0;
    else if( jump_type489_wr )
        jump_type489 <= wdata[31:0];
end


//jump_type490
assign jump_type490_reg[31:0]   = jump_type490                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type490 <= 32'h0;
    else if( jump_type490_wr )
        jump_type490 <= wdata[31:0];
end


//jump_type491
assign jump_type491_reg[31:0]   = jump_type491                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type491 <= 32'h0;
    else if( jump_type491_wr )
        jump_type491 <= wdata[31:0];
end


//jump_type492
assign jump_type492_reg[31:0]   = jump_type492                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type492 <= 32'h0;
    else if( jump_type492_wr )
        jump_type492 <= wdata[31:0];
end


//jump_type493
assign jump_type493_reg[31:0]   = jump_type493                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type493 <= 32'h0;
    else if( jump_type493_wr )
        jump_type493 <= wdata[31:0];
end


//jump_type494
assign jump_type494_reg[31:0]   = jump_type494                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type494 <= 32'h0;
    else if( jump_type494_wr )
        jump_type494 <= wdata[31:0];
end


//jump_type495
assign jump_type495_reg[31:0]   = jump_type495                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type495 <= 32'h0;
    else if( jump_type495_wr )
        jump_type495 <= wdata[31:0];
end


//jump_type496
assign jump_type496_reg[31:0]   = jump_type496                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type496 <= 32'h0;
    else if( jump_type496_wr )
        jump_type496 <= wdata[31:0];
end


//jump_type497
assign jump_type497_reg[31:0]   = jump_type497                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type497 <= 32'h0;
    else if( jump_type497_wr )
        jump_type497 <= wdata[31:0];
end


//jump_type498
assign jump_type498_reg[31:0]   = jump_type498                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type498 <= 32'h0;
    else if( jump_type498_wr )
        jump_type498 <= wdata[31:0];
end


//jump_type499
assign jump_type499_reg[31:0]   = jump_type499                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type499 <= 32'h0;
    else if( jump_type499_wr )
        jump_type499 <= wdata[31:0];
end


//jump_type500
assign jump_type500_reg[31:0]   = jump_type500                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type500 <= 32'h0;
    else if( jump_type500_wr )
        jump_type500 <= wdata[31:0];
end


//jump_type501
assign jump_type501_reg[31:0]   = jump_type501                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type501 <= 32'h0;
    else if( jump_type501_wr )
        jump_type501 <= wdata[31:0];
end


//jump_type502
assign jump_type502_reg[31:0]   = jump_type502                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type502 <= 32'h0;
    else if( jump_type502_wr )
        jump_type502 <= wdata[31:0];
end


//jump_type503
assign jump_type503_reg[31:0]   = jump_type503                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type503 <= 32'h0;
    else if( jump_type503_wr )
        jump_type503 <= wdata[31:0];
end


//jump_type504
assign jump_type504_reg[31:0]   = jump_type504                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type504 <= 32'h0;
    else if( jump_type504_wr )
        jump_type504 <= wdata[31:0];
end


//jump_type505
assign jump_type505_reg[31:0]   = jump_type505                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type505 <= 32'h0;
    else if( jump_type505_wr )
        jump_type505 <= wdata[31:0];
end


//jump_type506
assign jump_type506_reg[31:0]   = jump_type506                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type506 <= 32'h0;
    else if( jump_type506_wr )
        jump_type506 <= wdata[31:0];
end


//jump_type507
assign jump_type507_reg[31:0]   = jump_type507                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type507 <= 32'h0;
    else if( jump_type507_wr )
        jump_type507 <= wdata[31:0];
end


//jump_type508
assign jump_type508_reg[31:0]   = jump_type508                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type508 <= 32'h0;
    else if( jump_type508_wr )
        jump_type508 <= wdata[31:0];
end


//jump_type509
assign jump_type509_reg[31:0]   = jump_type509                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type509 <= 32'h0;
    else if( jump_type509_wr )
        jump_type509 <= wdata[31:0];
end


//jump_type510
assign jump_type510_reg[31:0]   = jump_type510                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type510 <= 32'h0;
    else if( jump_type510_wr )
        jump_type510 <= wdata[31:0];
end


//jump_type511
assign jump_type511_reg[31:28]  = 4'h0                        ;
assign jump_type511_reg[27:0]   = jump_type511                ;
always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        jump_type511 <= 28'h0;
    else if( jump_type511_wr )
        jump_type511 <= wdata[27:0];
end


//merger interrupt with group

//read
reg        [32-1:0]        rdata_tmp;
always @ ( * )
begin
    if ( ren )
    begin
        case( raddr )
            COMMON_PARA_REG:
                rdata_tmp = common_para_reg;
            JUMP_TYPE0_REG:
                rdata_tmp = jump_type0_reg;
            JUMP_TYPE1_REG:
                rdata_tmp = jump_type1_reg;
            JUMP_TYPE2_REG:
                rdata_tmp = jump_type2_reg;
            JUMP_TYPE3_REG:
                rdata_tmp = jump_type3_reg;
            JUMP_TYPE4_REG:
                rdata_tmp = jump_type4_reg;
            JUMP_TYPE5_REG:
                rdata_tmp = jump_type5_reg;
            JUMP_TYPE6_REG:
                rdata_tmp = jump_type6_reg;
            JUMP_TYPE7_REG:
                rdata_tmp = jump_type7_reg;
            JUMP_TYPE8_REG:
                rdata_tmp = jump_type8_reg;
            JUMP_TYPE9_REG:
                rdata_tmp = jump_type9_reg;
            JUMP_TYPE10_REG:
                rdata_tmp = jump_type10_reg;
            JUMP_TYPE11_REG:
                rdata_tmp = jump_type11_reg;
            JUMP_TYPE12_REG:
                rdata_tmp = jump_type12_reg;
            JUMP_TYPE13_REG:
                rdata_tmp = jump_type13_reg;
            JUMP_TYPE14_REG:
                rdata_tmp = jump_type14_reg;
            JUMP_TYPE15_REG:
                rdata_tmp = jump_type15_reg;
            JUMP_TYPE16_REG:
                rdata_tmp = jump_type16_reg;
            JUMP_TYPE17_REG:
                rdata_tmp = jump_type17_reg;
            JUMP_TYPE18_REG:
                rdata_tmp = jump_type18_reg;
            JUMP_TYPE19_REG:
                rdata_tmp = jump_type19_reg;
            JUMP_TYPE20_REG:
                rdata_tmp = jump_type20_reg;
            JUMP_TYPE21_REG:
                rdata_tmp = jump_type21_reg;
            JUMP_TYPE22_REG:
                rdata_tmp = jump_type22_reg;
            JUMP_TYPE23_REG:
                rdata_tmp = jump_type23_reg;
            JUMP_TYPE24_REG:
                rdata_tmp = jump_type24_reg;
            JUMP_TYPE25_REG:
                rdata_tmp = jump_type25_reg;
            JUMP_TYPE26_REG:
                rdata_tmp = jump_type26_reg;
            JUMP_TYPE27_REG:
                rdata_tmp = jump_type27_reg;
            JUMP_TYPE28_REG:
                rdata_tmp = jump_type28_reg;
            JUMP_TYPE29_REG:
                rdata_tmp = jump_type29_reg;
            JUMP_TYPE30_REG:
                rdata_tmp = jump_type30_reg;
            JUMP_TYPE31_REG:
                rdata_tmp = jump_type31_reg;
            JUMP_TYPE32_REG:
                rdata_tmp = jump_type32_reg;
            JUMP_TYPE33_REG:
                rdata_tmp = jump_type33_reg;
            JUMP_TYPE34_REG:
                rdata_tmp = jump_type34_reg;
            JUMP_TYPE35_REG:
                rdata_tmp = jump_type35_reg;
            JUMP_TYPE36_REG:
                rdata_tmp = jump_type36_reg;
            JUMP_TYPE37_REG:
                rdata_tmp = jump_type37_reg;
            JUMP_TYPE38_REG:
                rdata_tmp = jump_type38_reg;
            JUMP_TYPE39_REG:
                rdata_tmp = jump_type39_reg;
            JUMP_TYPE40_REG:
                rdata_tmp = jump_type40_reg;
            JUMP_TYPE41_REG:
                rdata_tmp = jump_type41_reg;
            JUMP_TYPE42_REG:
                rdata_tmp = jump_type42_reg;
            JUMP_TYPE43_REG:
                rdata_tmp = jump_type43_reg;
            JUMP_TYPE44_REG:
                rdata_tmp = jump_type44_reg;
            JUMP_TYPE45_REG:
                rdata_tmp = jump_type45_reg;
            JUMP_TYPE46_REG:
                rdata_tmp = jump_type46_reg;
            JUMP_TYPE47_REG:
                rdata_tmp = jump_type47_reg;
            JUMP_TYPE48_REG:
                rdata_tmp = jump_type48_reg;
            JUMP_TYPE49_REG:
                rdata_tmp = jump_type49_reg;
            JUMP_TYPE50_REG:
                rdata_tmp = jump_type50_reg;
            JUMP_TYPE51_REG:
                rdata_tmp = jump_type51_reg;
            JUMP_TYPE52_REG:
                rdata_tmp = jump_type52_reg;
            JUMP_TYPE53_REG:
                rdata_tmp = jump_type53_reg;
            JUMP_TYPE54_REG:
                rdata_tmp = jump_type54_reg;
            JUMP_TYPE55_REG:
                rdata_tmp = jump_type55_reg;
            JUMP_TYPE56_REG:
                rdata_tmp = jump_type56_reg;
            JUMP_TYPE57_REG:
                rdata_tmp = jump_type57_reg;
            JUMP_TYPE58_REG:
                rdata_tmp = jump_type58_reg;
            JUMP_TYPE59_REG:
                rdata_tmp = jump_type59_reg;
            JUMP_TYPE60_REG:
                rdata_tmp = jump_type60_reg;
            JUMP_TYPE61_REG:
                rdata_tmp = jump_type61_reg;
            JUMP_TYPE62_REG:
                rdata_tmp = jump_type62_reg;
            JUMP_TYPE63_REG:
                rdata_tmp = jump_type63_reg;
            JUMP_TYPE64_REG:
                rdata_tmp = jump_type64_reg;
            JUMP_TYPE65_REG:
                rdata_tmp = jump_type65_reg;
            JUMP_TYPE66_REG:
                rdata_tmp = jump_type66_reg;
            JUMP_TYPE67_REG:
                rdata_tmp = jump_type67_reg;
            JUMP_TYPE68_REG:
                rdata_tmp = jump_type68_reg;
            JUMP_TYPE69_REG:
                rdata_tmp = jump_type69_reg;
            JUMP_TYPE70_REG:
                rdata_tmp = jump_type70_reg;
            JUMP_TYPE71_REG:
                rdata_tmp = jump_type71_reg;
            JUMP_TYPE72_REG:
                rdata_tmp = jump_type72_reg;
            JUMP_TYPE73_REG:
                rdata_tmp = jump_type73_reg;
            JUMP_TYPE74_REG:
                rdata_tmp = jump_type74_reg;
            JUMP_TYPE75_REG:
                rdata_tmp = jump_type75_reg;
            JUMP_TYPE76_REG:
                rdata_tmp = jump_type76_reg;
            JUMP_TYPE77_REG:
                rdata_tmp = jump_type77_reg;
            JUMP_TYPE78_REG:
                rdata_tmp = jump_type78_reg;
            JUMP_TYPE79_REG:
                rdata_tmp = jump_type79_reg;
            JUMP_TYPE80_REG:
                rdata_tmp = jump_type80_reg;
            JUMP_TYPE81_REG:
                rdata_tmp = jump_type81_reg;
            JUMP_TYPE82_REG:
                rdata_tmp = jump_type82_reg;
            JUMP_TYPE83_REG:
                rdata_tmp = jump_type83_reg;
            JUMP_TYPE84_REG:
                rdata_tmp = jump_type84_reg;
            JUMP_TYPE85_REG:
                rdata_tmp = jump_type85_reg;
            JUMP_TYPE86_REG:
                rdata_tmp = jump_type86_reg;
            JUMP_TYPE87_REG:
                rdata_tmp = jump_type87_reg;
            JUMP_TYPE88_REG:
                rdata_tmp = jump_type88_reg;
            JUMP_TYPE89_REG:
                rdata_tmp = jump_type89_reg;
            JUMP_TYPE90_REG:
                rdata_tmp = jump_type90_reg;
            JUMP_TYPE91_REG:
                rdata_tmp = jump_type91_reg;
            JUMP_TYPE92_REG:
                rdata_tmp = jump_type92_reg;
            JUMP_TYPE93_REG:
                rdata_tmp = jump_type93_reg;
            JUMP_TYPE94_REG:
                rdata_tmp = jump_type94_reg;
            JUMP_TYPE95_REG:
                rdata_tmp = jump_type95_reg;
            JUMP_TYPE96_REG:
                rdata_tmp = jump_type96_reg;
            JUMP_TYPE97_REG:
                rdata_tmp = jump_type97_reg;
            JUMP_TYPE98_REG:
                rdata_tmp = jump_type98_reg;
            JUMP_TYPE99_REG:
                rdata_tmp = jump_type99_reg;
            JUMP_TYPE100_REG:
                rdata_tmp = jump_type100_reg;
            JUMP_TYPE101_REG:
                rdata_tmp = jump_type101_reg;
            JUMP_TYPE102_REG:
                rdata_tmp = jump_type102_reg;
            JUMP_TYPE103_REG:
                rdata_tmp = jump_type103_reg;
            JUMP_TYPE104_REG:
                rdata_tmp = jump_type104_reg;
            JUMP_TYPE105_REG:
                rdata_tmp = jump_type105_reg;
            JUMP_TYPE106_REG:
                rdata_tmp = jump_type106_reg;
            JUMP_TYPE107_REG:
                rdata_tmp = jump_type107_reg;
            JUMP_TYPE108_REG:
                rdata_tmp = jump_type108_reg;
            JUMP_TYPE109_REG:
                rdata_tmp = jump_type109_reg;
            JUMP_TYPE110_REG:
                rdata_tmp = jump_type110_reg;
            JUMP_TYPE111_REG:
                rdata_tmp = jump_type111_reg;
            JUMP_TYPE112_REG:
                rdata_tmp = jump_type112_reg;
            JUMP_TYPE113_REG:
                rdata_tmp = jump_type113_reg;
            JUMP_TYPE114_REG:
                rdata_tmp = jump_type114_reg;
            JUMP_TYPE115_REG:
                rdata_tmp = jump_type115_reg;
            JUMP_TYPE116_REG:
                rdata_tmp = jump_type116_reg;
            JUMP_TYPE117_REG:
                rdata_tmp = jump_type117_reg;
            JUMP_TYPE118_REG:
                rdata_tmp = jump_type118_reg;
            JUMP_TYPE119_REG:
                rdata_tmp = jump_type119_reg;
            JUMP_TYPE120_REG:
                rdata_tmp = jump_type120_reg;
            JUMP_TYPE121_REG:
                rdata_tmp = jump_type121_reg;
            JUMP_TYPE122_REG:
                rdata_tmp = jump_type122_reg;
            JUMP_TYPE123_REG:
                rdata_tmp = jump_type123_reg;
            JUMP_TYPE124_REG:
                rdata_tmp = jump_type124_reg;
            JUMP_TYPE125_REG:
                rdata_tmp = jump_type125_reg;
            JUMP_TYPE126_REG:
                rdata_tmp = jump_type126_reg;
            JUMP_TYPE127_REG:
                rdata_tmp = jump_type127_reg;
            JUMP_TYPE128_REG:
                rdata_tmp = jump_type128_reg;
            JUMP_TYPE129_REG:
                rdata_tmp = jump_type129_reg;
            JUMP_TYPE130_REG:
                rdata_tmp = jump_type130_reg;
            JUMP_TYPE131_REG:
                rdata_tmp = jump_type131_reg;
            JUMP_TYPE132_REG:
                rdata_tmp = jump_type132_reg;
            JUMP_TYPE133_REG:
                rdata_tmp = jump_type133_reg;
            JUMP_TYPE134_REG:
                rdata_tmp = jump_type134_reg;
            JUMP_TYPE135_REG:
                rdata_tmp = jump_type135_reg;
            JUMP_TYPE136_REG:
                rdata_tmp = jump_type136_reg;
            JUMP_TYPE137_REG:
                rdata_tmp = jump_type137_reg;
            JUMP_TYPE138_REG:
                rdata_tmp = jump_type138_reg;
            JUMP_TYPE139_REG:
                rdata_tmp = jump_type139_reg;
            JUMP_TYPE140_REG:
                rdata_tmp = jump_type140_reg;
            JUMP_TYPE141_REG:
                rdata_tmp = jump_type141_reg;
            JUMP_TYPE142_REG:
                rdata_tmp = jump_type142_reg;
            JUMP_TYPE143_REG:
                rdata_tmp = jump_type143_reg;
            JUMP_TYPE144_REG:
                rdata_tmp = jump_type144_reg;
            JUMP_TYPE145_REG:
                rdata_tmp = jump_type145_reg;
            JUMP_TYPE146_REG:
                rdata_tmp = jump_type146_reg;
            JUMP_TYPE147_REG:
                rdata_tmp = jump_type147_reg;
            JUMP_TYPE148_REG:
                rdata_tmp = jump_type148_reg;
            JUMP_TYPE149_REG:
                rdata_tmp = jump_type149_reg;
            JUMP_TYPE150_REG:
                rdata_tmp = jump_type150_reg;
            JUMP_TYPE151_REG:
                rdata_tmp = jump_type151_reg;
            JUMP_TYPE152_REG:
                rdata_tmp = jump_type152_reg;
            JUMP_TYPE153_REG:
                rdata_tmp = jump_type153_reg;
            JUMP_TYPE154_REG:
                rdata_tmp = jump_type154_reg;
            JUMP_TYPE155_REG:
                rdata_tmp = jump_type155_reg;
            JUMP_TYPE156_REG:
                rdata_tmp = jump_type156_reg;
            JUMP_TYPE157_REG:
                rdata_tmp = jump_type157_reg;
            JUMP_TYPE158_REG:
                rdata_tmp = jump_type158_reg;
            JUMP_TYPE159_REG:
                rdata_tmp = jump_type159_reg;
            JUMP_TYPE160_REG:
                rdata_tmp = jump_type160_reg;
            JUMP_TYPE161_REG:
                rdata_tmp = jump_type161_reg;
            JUMP_TYPE162_REG:
                rdata_tmp = jump_type162_reg;
            JUMP_TYPE163_REG:
                rdata_tmp = jump_type163_reg;
            JUMP_TYPE164_REG:
                rdata_tmp = jump_type164_reg;
            JUMP_TYPE165_REG:
                rdata_tmp = jump_type165_reg;
            JUMP_TYPE166_REG:
                rdata_tmp = jump_type166_reg;
            JUMP_TYPE167_REG:
                rdata_tmp = jump_type167_reg;
            JUMP_TYPE168_REG:
                rdata_tmp = jump_type168_reg;
            JUMP_TYPE169_REG:
                rdata_tmp = jump_type169_reg;
            JUMP_TYPE170_REG:
                rdata_tmp = jump_type170_reg;
            JUMP_TYPE171_REG:
                rdata_tmp = jump_type171_reg;
            JUMP_TYPE172_REG:
                rdata_tmp = jump_type172_reg;
            JUMP_TYPE173_REG:
                rdata_tmp = jump_type173_reg;
            JUMP_TYPE174_REG:
                rdata_tmp = jump_type174_reg;
            JUMP_TYPE175_REG:
                rdata_tmp = jump_type175_reg;
            JUMP_TYPE176_REG:
                rdata_tmp = jump_type176_reg;
            JUMP_TYPE177_REG:
                rdata_tmp = jump_type177_reg;
            JUMP_TYPE178_REG:
                rdata_tmp = jump_type178_reg;
            JUMP_TYPE179_REG:
                rdata_tmp = jump_type179_reg;
            JUMP_TYPE180_REG:
                rdata_tmp = jump_type180_reg;
            JUMP_TYPE181_REG:
                rdata_tmp = jump_type181_reg;
            JUMP_TYPE182_REG:
                rdata_tmp = jump_type182_reg;
            JUMP_TYPE183_REG:
                rdata_tmp = jump_type183_reg;
            JUMP_TYPE184_REG:
                rdata_tmp = jump_type184_reg;
            JUMP_TYPE185_REG:
                rdata_tmp = jump_type185_reg;
            JUMP_TYPE186_REG:
                rdata_tmp = jump_type186_reg;
            JUMP_TYPE187_REG:
                rdata_tmp = jump_type187_reg;
            JUMP_TYPE188_REG:
                rdata_tmp = jump_type188_reg;
            JUMP_TYPE189_REG:
                rdata_tmp = jump_type189_reg;
            JUMP_TYPE190_REG:
                rdata_tmp = jump_type190_reg;
            JUMP_TYPE191_REG:
                rdata_tmp = jump_type191_reg;
            JUMP_TYPE192_REG:
                rdata_tmp = jump_type192_reg;
            JUMP_TYPE193_REG:
                rdata_tmp = jump_type193_reg;
            JUMP_TYPE194_REG:
                rdata_tmp = jump_type194_reg;
            JUMP_TYPE195_REG:
                rdata_tmp = jump_type195_reg;
            JUMP_TYPE196_REG:
                rdata_tmp = jump_type196_reg;
            JUMP_TYPE197_REG:
                rdata_tmp = jump_type197_reg;
            JUMP_TYPE198_REG:
                rdata_tmp = jump_type198_reg;
            JUMP_TYPE199_REG:
                rdata_tmp = jump_type199_reg;
            JUMP_TYPE200_REG:
                rdata_tmp = jump_type200_reg;
            JUMP_TYPE201_REG:
                rdata_tmp = jump_type201_reg;
            JUMP_TYPE202_REG:
                rdata_tmp = jump_type202_reg;
            JUMP_TYPE203_REG:
                rdata_tmp = jump_type203_reg;
            JUMP_TYPE204_REG:
                rdata_tmp = jump_type204_reg;
            JUMP_TYPE205_REG:
                rdata_tmp = jump_type205_reg;
            JUMP_TYPE206_REG:
                rdata_tmp = jump_type206_reg;
            JUMP_TYPE207_REG:
                rdata_tmp = jump_type207_reg;
            JUMP_TYPE208_REG:
                rdata_tmp = jump_type208_reg;
            JUMP_TYPE209_REG:
                rdata_tmp = jump_type209_reg;
            JUMP_TYPE210_REG:
                rdata_tmp = jump_type210_reg;
            JUMP_TYPE211_REG:
                rdata_tmp = jump_type211_reg;
            JUMP_TYPE212_REG:
                rdata_tmp = jump_type212_reg;
            JUMP_TYPE213_REG:
                rdata_tmp = jump_type213_reg;
            JUMP_TYPE214_REG:
                rdata_tmp = jump_type214_reg;
            JUMP_TYPE215_REG:
                rdata_tmp = jump_type215_reg;
            JUMP_TYPE216_REG:
                rdata_tmp = jump_type216_reg;
            JUMP_TYPE217_REG:
                rdata_tmp = jump_type217_reg;
            JUMP_TYPE218_REG:
                rdata_tmp = jump_type218_reg;
            JUMP_TYPE219_REG:
                rdata_tmp = jump_type219_reg;
            JUMP_TYPE220_REG:
                rdata_tmp = jump_type220_reg;
            JUMP_TYPE221_REG:
                rdata_tmp = jump_type221_reg;
            JUMP_TYPE222_REG:
                rdata_tmp = jump_type222_reg;
            JUMP_TYPE223_REG:
                rdata_tmp = jump_type223_reg;
            JUMP_TYPE224_REG:
                rdata_tmp = jump_type224_reg;
            JUMP_TYPE225_REG:
                rdata_tmp = jump_type225_reg;
            JUMP_TYPE226_REG:
                rdata_tmp = jump_type226_reg;
            JUMP_TYPE227_REG:
                rdata_tmp = jump_type227_reg;
            JUMP_TYPE228_REG:
                rdata_tmp = jump_type228_reg;
            JUMP_TYPE229_REG:
                rdata_tmp = jump_type229_reg;
            JUMP_TYPE230_REG:
                rdata_tmp = jump_type230_reg;
            JUMP_TYPE231_REG:
                rdata_tmp = jump_type231_reg;
            JUMP_TYPE232_REG:
                rdata_tmp = jump_type232_reg;
            JUMP_TYPE233_REG:
                rdata_tmp = jump_type233_reg;
            JUMP_TYPE234_REG:
                rdata_tmp = jump_type234_reg;
            JUMP_TYPE235_REG:
                rdata_tmp = jump_type235_reg;
            JUMP_TYPE236_REG:
                rdata_tmp = jump_type236_reg;
            JUMP_TYPE237_REG:
                rdata_tmp = jump_type237_reg;
            JUMP_TYPE238_REG:
                rdata_tmp = jump_type238_reg;
            JUMP_TYPE239_REG:
                rdata_tmp = jump_type239_reg;
            JUMP_TYPE240_REG:
                rdata_tmp = jump_type240_reg;
            JUMP_TYPE241_REG:
                rdata_tmp = jump_type241_reg;
            JUMP_TYPE242_REG:
                rdata_tmp = jump_type242_reg;
            JUMP_TYPE243_REG:
                rdata_tmp = jump_type243_reg;
            JUMP_TYPE244_REG:
                rdata_tmp = jump_type244_reg;
            JUMP_TYPE245_REG:
                rdata_tmp = jump_type245_reg;
            JUMP_TYPE246_REG:
                rdata_tmp = jump_type246_reg;
            JUMP_TYPE247_REG:
                rdata_tmp = jump_type247_reg;
            JUMP_TYPE248_REG:
                rdata_tmp = jump_type248_reg;
            JUMP_TYPE249_REG:
                rdata_tmp = jump_type249_reg;
            JUMP_TYPE250_REG:
                rdata_tmp = jump_type250_reg;
            JUMP_TYPE251_REG:
                rdata_tmp = jump_type251_reg;
            JUMP_TYPE252_REG:
                rdata_tmp = jump_type252_reg;
            JUMP_TYPE253_REG:
                rdata_tmp = jump_type253_reg;
            JUMP_TYPE254_REG:
                rdata_tmp = jump_type254_reg;
            JUMP_TYPE255_REG:
                rdata_tmp = jump_type255_reg;
            JUMP_TYPE256_REG:
                rdata_tmp = jump_type256_reg;
            JUMP_TYPE257_REG:
                rdata_tmp = jump_type257_reg;
            JUMP_TYPE258_REG:
                rdata_tmp = jump_type258_reg;
            JUMP_TYPE259_REG:
                rdata_tmp = jump_type259_reg;
            JUMP_TYPE260_REG:
                rdata_tmp = jump_type260_reg;
            JUMP_TYPE261_REG:
                rdata_tmp = jump_type261_reg;
            JUMP_TYPE262_REG:
                rdata_tmp = jump_type262_reg;
            JUMP_TYPE263_REG:
                rdata_tmp = jump_type263_reg;
            JUMP_TYPE264_REG:
                rdata_tmp = jump_type264_reg;
            JUMP_TYPE265_REG:
                rdata_tmp = jump_type265_reg;
            JUMP_TYPE266_REG:
                rdata_tmp = jump_type266_reg;
            JUMP_TYPE267_REG:
                rdata_tmp = jump_type267_reg;
            JUMP_TYPE268_REG:
                rdata_tmp = jump_type268_reg;
            JUMP_TYPE269_REG:
                rdata_tmp = jump_type269_reg;
            JUMP_TYPE270_REG:
                rdata_tmp = jump_type270_reg;
            JUMP_TYPE271_REG:
                rdata_tmp = jump_type271_reg;
            JUMP_TYPE272_REG:
                rdata_tmp = jump_type272_reg;
            JUMP_TYPE273_REG:
                rdata_tmp = jump_type273_reg;
            JUMP_TYPE274_REG:
                rdata_tmp = jump_type274_reg;
            JUMP_TYPE275_REG:
                rdata_tmp = jump_type275_reg;
            JUMP_TYPE276_REG:
                rdata_tmp = jump_type276_reg;
            JUMP_TYPE277_REG:
                rdata_tmp = jump_type277_reg;
            JUMP_TYPE278_REG:
                rdata_tmp = jump_type278_reg;
            JUMP_TYPE279_REG:
                rdata_tmp = jump_type279_reg;
            JUMP_TYPE280_REG:
                rdata_tmp = jump_type280_reg;
            JUMP_TYPE281_REG:
                rdata_tmp = jump_type281_reg;
            JUMP_TYPE282_REG:
                rdata_tmp = jump_type282_reg;
            JUMP_TYPE283_REG:
                rdata_tmp = jump_type283_reg;
            JUMP_TYPE284_REG:
                rdata_tmp = jump_type284_reg;
            JUMP_TYPE285_REG:
                rdata_tmp = jump_type285_reg;
            JUMP_TYPE286_REG:
                rdata_tmp = jump_type286_reg;
            JUMP_TYPE287_REG:
                rdata_tmp = jump_type287_reg;
            JUMP_TYPE288_REG:
                rdata_tmp = jump_type288_reg;
            JUMP_TYPE289_REG:
                rdata_tmp = jump_type289_reg;
            JUMP_TYPE290_REG:
                rdata_tmp = jump_type290_reg;
            JUMP_TYPE291_REG:
                rdata_tmp = jump_type291_reg;
            JUMP_TYPE292_REG:
                rdata_tmp = jump_type292_reg;
            JUMP_TYPE293_REG:
                rdata_tmp = jump_type293_reg;
            JUMP_TYPE294_REG:
                rdata_tmp = jump_type294_reg;
            JUMP_TYPE295_REG:
                rdata_tmp = jump_type295_reg;
            JUMP_TYPE296_REG:
                rdata_tmp = jump_type296_reg;
            JUMP_TYPE297_REG:
                rdata_tmp = jump_type297_reg;
            JUMP_TYPE298_REG:
                rdata_tmp = jump_type298_reg;
            JUMP_TYPE299_REG:
                rdata_tmp = jump_type299_reg;
            JUMP_TYPE300_REG:
                rdata_tmp = jump_type300_reg;
            JUMP_TYPE301_REG:
                rdata_tmp = jump_type301_reg;
            JUMP_TYPE302_REG:
                rdata_tmp = jump_type302_reg;
            JUMP_TYPE303_REG:
                rdata_tmp = jump_type303_reg;
            JUMP_TYPE304_REG:
                rdata_tmp = jump_type304_reg;
            JUMP_TYPE305_REG:
                rdata_tmp = jump_type305_reg;
            JUMP_TYPE306_REG:
                rdata_tmp = jump_type306_reg;
            JUMP_TYPE307_REG:
                rdata_tmp = jump_type307_reg;
            JUMP_TYPE308_REG:
                rdata_tmp = jump_type308_reg;
            JUMP_TYPE309_REG:
                rdata_tmp = jump_type309_reg;
            JUMP_TYPE310_REG:
                rdata_tmp = jump_type310_reg;
            JUMP_TYPE311_REG:
                rdata_tmp = jump_type311_reg;
            JUMP_TYPE312_REG:
                rdata_tmp = jump_type312_reg;
            JUMP_TYPE313_REG:
                rdata_tmp = jump_type313_reg;
            JUMP_TYPE314_REG:
                rdata_tmp = jump_type314_reg;
            JUMP_TYPE315_REG:
                rdata_tmp = jump_type315_reg;
            JUMP_TYPE316_REG:
                rdata_tmp = jump_type316_reg;
            JUMP_TYPE317_REG:
                rdata_tmp = jump_type317_reg;
            JUMP_TYPE318_REG:
                rdata_tmp = jump_type318_reg;
            JUMP_TYPE319_REG:
                rdata_tmp = jump_type319_reg;
            JUMP_TYPE320_REG:
                rdata_tmp = jump_type320_reg;
            JUMP_TYPE321_REG:
                rdata_tmp = jump_type321_reg;
            JUMP_TYPE322_REG:
                rdata_tmp = jump_type322_reg;
            JUMP_TYPE323_REG:
                rdata_tmp = jump_type323_reg;
            JUMP_TYPE324_REG:
                rdata_tmp = jump_type324_reg;
            JUMP_TYPE325_REG:
                rdata_tmp = jump_type325_reg;
            JUMP_TYPE326_REG:
                rdata_tmp = jump_type326_reg;
            JUMP_TYPE327_REG:
                rdata_tmp = jump_type327_reg;
            JUMP_TYPE328_REG:
                rdata_tmp = jump_type328_reg;
            JUMP_TYPE329_REG:
                rdata_tmp = jump_type329_reg;
            JUMP_TYPE330_REG:
                rdata_tmp = jump_type330_reg;
            JUMP_TYPE331_REG:
                rdata_tmp = jump_type331_reg;
            JUMP_TYPE332_REG:
                rdata_tmp = jump_type332_reg;
            JUMP_TYPE333_REG:
                rdata_tmp = jump_type333_reg;
            JUMP_TYPE334_REG:
                rdata_tmp = jump_type334_reg;
            JUMP_TYPE335_REG:
                rdata_tmp = jump_type335_reg;
            JUMP_TYPE336_REG:
                rdata_tmp = jump_type336_reg;
            JUMP_TYPE337_REG:
                rdata_tmp = jump_type337_reg;
            JUMP_TYPE338_REG:
                rdata_tmp = jump_type338_reg;
            JUMP_TYPE339_REG:
                rdata_tmp = jump_type339_reg;
            JUMP_TYPE340_REG:
                rdata_tmp = jump_type340_reg;
            JUMP_TYPE341_REG:
                rdata_tmp = jump_type341_reg;
            JUMP_TYPE342_REG:
                rdata_tmp = jump_type342_reg;
            JUMP_TYPE343_REG:
                rdata_tmp = jump_type343_reg;
            JUMP_TYPE344_REG:
                rdata_tmp = jump_type344_reg;
            JUMP_TYPE345_REG:
                rdata_tmp = jump_type345_reg;
            JUMP_TYPE346_REG:
                rdata_tmp = jump_type346_reg;
            JUMP_TYPE347_REG:
                rdata_tmp = jump_type347_reg;
            JUMP_TYPE348_REG:
                rdata_tmp = jump_type348_reg;
            JUMP_TYPE349_REG:
                rdata_tmp = jump_type349_reg;
            JUMP_TYPE350_REG:
                rdata_tmp = jump_type350_reg;
            JUMP_TYPE351_REG:
                rdata_tmp = jump_type351_reg;
            JUMP_TYPE352_REG:
                rdata_tmp = jump_type352_reg;
            JUMP_TYPE353_REG:
                rdata_tmp = jump_type353_reg;
            JUMP_TYPE354_REG:
                rdata_tmp = jump_type354_reg;
            JUMP_TYPE355_REG:
                rdata_tmp = jump_type355_reg;
            JUMP_TYPE356_REG:
                rdata_tmp = jump_type356_reg;
            JUMP_TYPE357_REG:
                rdata_tmp = jump_type357_reg;
            JUMP_TYPE358_REG:
                rdata_tmp = jump_type358_reg;
            JUMP_TYPE359_REG:
                rdata_tmp = jump_type359_reg;
            JUMP_TYPE360_REG:
                rdata_tmp = jump_type360_reg;
            JUMP_TYPE361_REG:
                rdata_tmp = jump_type361_reg;
            JUMP_TYPE362_REG:
                rdata_tmp = jump_type362_reg;
            JUMP_TYPE363_REG:
                rdata_tmp = jump_type363_reg;
            JUMP_TYPE364_REG:
                rdata_tmp = jump_type364_reg;
            JUMP_TYPE365_REG:
                rdata_tmp = jump_type365_reg;
            JUMP_TYPE366_REG:
                rdata_tmp = jump_type366_reg;
            JUMP_TYPE367_REG:
                rdata_tmp = jump_type367_reg;
            JUMP_TYPE368_REG:
                rdata_tmp = jump_type368_reg;
            JUMP_TYPE369_REG:
                rdata_tmp = jump_type369_reg;
            JUMP_TYPE370_REG:
                rdata_tmp = jump_type370_reg;
            JUMP_TYPE371_REG:
                rdata_tmp = jump_type371_reg;
            JUMP_TYPE372_REG:
                rdata_tmp = jump_type372_reg;
            JUMP_TYPE373_REG:
                rdata_tmp = jump_type373_reg;
            JUMP_TYPE374_REG:
                rdata_tmp = jump_type374_reg;
            JUMP_TYPE375_REG:
                rdata_tmp = jump_type375_reg;
            JUMP_TYPE376_REG:
                rdata_tmp = jump_type376_reg;
            JUMP_TYPE377_REG:
                rdata_tmp = jump_type377_reg;
            JUMP_TYPE378_REG:
                rdata_tmp = jump_type378_reg;
            JUMP_TYPE379_REG:
                rdata_tmp = jump_type379_reg;
            JUMP_TYPE380_REG:
                rdata_tmp = jump_type380_reg;
            JUMP_TYPE381_REG:
                rdata_tmp = jump_type381_reg;
            JUMP_TYPE382_REG:
                rdata_tmp = jump_type382_reg;
            JUMP_TYPE383_REG:
                rdata_tmp = jump_type383_reg;
            JUMP_TYPE384_REG:
                rdata_tmp = jump_type384_reg;
            JUMP_TYPE385_REG:
                rdata_tmp = jump_type385_reg;
            JUMP_TYPE386_REG:
                rdata_tmp = jump_type386_reg;
            JUMP_TYPE387_REG:
                rdata_tmp = jump_type387_reg;
            JUMP_TYPE388_REG:
                rdata_tmp = jump_type388_reg;
            JUMP_TYPE389_REG:
                rdata_tmp = jump_type389_reg;
            JUMP_TYPE390_REG:
                rdata_tmp = jump_type390_reg;
            JUMP_TYPE391_REG:
                rdata_tmp = jump_type391_reg;
            JUMP_TYPE392_REG:
                rdata_tmp = jump_type392_reg;
            JUMP_TYPE393_REG:
                rdata_tmp = jump_type393_reg;
            JUMP_TYPE394_REG:
                rdata_tmp = jump_type394_reg;
            JUMP_TYPE395_REG:
                rdata_tmp = jump_type395_reg;
            JUMP_TYPE396_REG:
                rdata_tmp = jump_type396_reg;
            JUMP_TYPE397_REG:
                rdata_tmp = jump_type397_reg;
            JUMP_TYPE398_REG:
                rdata_tmp = jump_type398_reg;
            JUMP_TYPE399_REG:
                rdata_tmp = jump_type399_reg;
            JUMP_TYPE400_REG:
                rdata_tmp = jump_type400_reg;
            JUMP_TYPE401_REG:
                rdata_tmp = jump_type401_reg;
            JUMP_TYPE402_REG:
                rdata_tmp = jump_type402_reg;
            JUMP_TYPE403_REG:
                rdata_tmp = jump_type403_reg;
            JUMP_TYPE404_REG:
                rdata_tmp = jump_type404_reg;
            JUMP_TYPE405_REG:
                rdata_tmp = jump_type405_reg;
            JUMP_TYPE406_REG:
                rdata_tmp = jump_type406_reg;
            JUMP_TYPE407_REG:
                rdata_tmp = jump_type407_reg;
            JUMP_TYPE408_REG:
                rdata_tmp = jump_type408_reg;
            JUMP_TYPE409_REG:
                rdata_tmp = jump_type409_reg;
            JUMP_TYPE410_REG:
                rdata_tmp = jump_type410_reg;
            JUMP_TYPE411_REG:
                rdata_tmp = jump_type411_reg;
            JUMP_TYPE412_REG:
                rdata_tmp = jump_type412_reg;
            JUMP_TYPE413_REG:
                rdata_tmp = jump_type413_reg;
            JUMP_TYPE414_REG:
                rdata_tmp = jump_type414_reg;
            JUMP_TYPE415_REG:
                rdata_tmp = jump_type415_reg;
            JUMP_TYPE416_REG:
                rdata_tmp = jump_type416_reg;
            JUMP_TYPE417_REG:
                rdata_tmp = jump_type417_reg;
            JUMP_TYPE418_REG:
                rdata_tmp = jump_type418_reg;
            JUMP_TYPE419_REG:
                rdata_tmp = jump_type419_reg;
            JUMP_TYPE420_REG:
                rdata_tmp = jump_type420_reg;
            JUMP_TYPE421_REG:
                rdata_tmp = jump_type421_reg;
            JUMP_TYPE422_REG:
                rdata_tmp = jump_type422_reg;
            JUMP_TYPE423_REG:
                rdata_tmp = jump_type423_reg;
            JUMP_TYPE424_REG:
                rdata_tmp = jump_type424_reg;
            JUMP_TYPE425_REG:
                rdata_tmp = jump_type425_reg;
            JUMP_TYPE426_REG:
                rdata_tmp = jump_type426_reg;
            JUMP_TYPE427_REG:
                rdata_tmp = jump_type427_reg;
            JUMP_TYPE428_REG:
                rdata_tmp = jump_type428_reg;
            JUMP_TYPE429_REG:
                rdata_tmp = jump_type429_reg;
            JUMP_TYPE430_REG:
                rdata_tmp = jump_type430_reg;
            JUMP_TYPE431_REG:
                rdata_tmp = jump_type431_reg;
            JUMP_TYPE432_REG:
                rdata_tmp = jump_type432_reg;
            JUMP_TYPE433_REG:
                rdata_tmp = jump_type433_reg;
            JUMP_TYPE434_REG:
                rdata_tmp = jump_type434_reg;
            JUMP_TYPE435_REG:
                rdata_tmp = jump_type435_reg;
            JUMP_TYPE436_REG:
                rdata_tmp = jump_type436_reg;
            JUMP_TYPE437_REG:
                rdata_tmp = jump_type437_reg;
            JUMP_TYPE438_REG:
                rdata_tmp = jump_type438_reg;
            JUMP_TYPE439_REG:
                rdata_tmp = jump_type439_reg;
            JUMP_TYPE440_REG:
                rdata_tmp = jump_type440_reg;
            JUMP_TYPE441_REG:
                rdata_tmp = jump_type441_reg;
            JUMP_TYPE442_REG:
                rdata_tmp = jump_type442_reg;
            JUMP_TYPE443_REG:
                rdata_tmp = jump_type443_reg;
            JUMP_TYPE444_REG:
                rdata_tmp = jump_type444_reg;
            JUMP_TYPE445_REG:
                rdata_tmp = jump_type445_reg;
            JUMP_TYPE446_REG:
                rdata_tmp = jump_type446_reg;
            JUMP_TYPE447_REG:
                rdata_tmp = jump_type447_reg;
            JUMP_TYPE448_REG:
                rdata_tmp = jump_type448_reg;
            JUMP_TYPE449_REG:
                rdata_tmp = jump_type449_reg;
            JUMP_TYPE450_REG:
                rdata_tmp = jump_type450_reg;
            JUMP_TYPE451_REG:
                rdata_tmp = jump_type451_reg;
            JUMP_TYPE452_REG:
                rdata_tmp = jump_type452_reg;
            JUMP_TYPE453_REG:
                rdata_tmp = jump_type453_reg;
            JUMP_TYPE454_REG:
                rdata_tmp = jump_type454_reg;
            JUMP_TYPE455_REG:
                rdata_tmp = jump_type455_reg;
            JUMP_TYPE456_REG:
                rdata_tmp = jump_type456_reg;
            JUMP_TYPE457_REG:
                rdata_tmp = jump_type457_reg;
            JUMP_TYPE458_REG:
                rdata_tmp = jump_type458_reg;
            JUMP_TYPE459_REG:
                rdata_tmp = jump_type459_reg;
            JUMP_TYPE460_REG:
                rdata_tmp = jump_type460_reg;
            JUMP_TYPE461_REG:
                rdata_tmp = jump_type461_reg;
            JUMP_TYPE462_REG:
                rdata_tmp = jump_type462_reg;
            JUMP_TYPE463_REG:
                rdata_tmp = jump_type463_reg;
            JUMP_TYPE464_REG:
                rdata_tmp = jump_type464_reg;
            JUMP_TYPE465_REG:
                rdata_tmp = jump_type465_reg;
            JUMP_TYPE466_REG:
                rdata_tmp = jump_type466_reg;
            JUMP_TYPE467_REG:
                rdata_tmp = jump_type467_reg;
            JUMP_TYPE468_REG:
                rdata_tmp = jump_type468_reg;
            JUMP_TYPE469_REG:
                rdata_tmp = jump_type469_reg;
            JUMP_TYPE470_REG:
                rdata_tmp = jump_type470_reg;
            JUMP_TYPE471_REG:
                rdata_tmp = jump_type471_reg;
            JUMP_TYPE472_REG:
                rdata_tmp = jump_type472_reg;
            JUMP_TYPE473_REG:
                rdata_tmp = jump_type473_reg;
            JUMP_TYPE474_REG:
                rdata_tmp = jump_type474_reg;
            JUMP_TYPE475_REG:
                rdata_tmp = jump_type475_reg;
            JUMP_TYPE476_REG:
                rdata_tmp = jump_type476_reg;
            JUMP_TYPE477_REG:
                rdata_tmp = jump_type477_reg;
            JUMP_TYPE478_REG:
                rdata_tmp = jump_type478_reg;
            JUMP_TYPE479_REG:
                rdata_tmp = jump_type479_reg;
            JUMP_TYPE480_REG:
                rdata_tmp = jump_type480_reg;
            JUMP_TYPE481_REG:
                rdata_tmp = jump_type481_reg;
            JUMP_TYPE482_REG:
                rdata_tmp = jump_type482_reg;
            JUMP_TYPE483_REG:
                rdata_tmp = jump_type483_reg;
            JUMP_TYPE484_REG:
                rdata_tmp = jump_type484_reg;
            JUMP_TYPE485_REG:
                rdata_tmp = jump_type485_reg;
            JUMP_TYPE486_REG:
                rdata_tmp = jump_type486_reg;
            JUMP_TYPE487_REG:
                rdata_tmp = jump_type487_reg;
            JUMP_TYPE488_REG:
                rdata_tmp = jump_type488_reg;
            JUMP_TYPE489_REG:
                rdata_tmp = jump_type489_reg;
            JUMP_TYPE490_REG:
                rdata_tmp = jump_type490_reg;
            JUMP_TYPE491_REG:
                rdata_tmp = jump_type491_reg;
            JUMP_TYPE492_REG:
                rdata_tmp = jump_type492_reg;
            JUMP_TYPE493_REG:
                rdata_tmp = jump_type493_reg;
            JUMP_TYPE494_REG:
                rdata_tmp = jump_type494_reg;
            JUMP_TYPE495_REG:
                rdata_tmp = jump_type495_reg;
            JUMP_TYPE496_REG:
                rdata_tmp = jump_type496_reg;
            JUMP_TYPE497_REG:
                rdata_tmp = jump_type497_reg;
            JUMP_TYPE498_REG:
                rdata_tmp = jump_type498_reg;
            JUMP_TYPE499_REG:
                rdata_tmp = jump_type499_reg;
            JUMP_TYPE500_REG:
                rdata_tmp = jump_type500_reg;
            JUMP_TYPE501_REG:
                rdata_tmp = jump_type501_reg;
            JUMP_TYPE502_REG:
                rdata_tmp = jump_type502_reg;
            JUMP_TYPE503_REG:
                rdata_tmp = jump_type503_reg;
            JUMP_TYPE504_REG:
                rdata_tmp = jump_type504_reg;
            JUMP_TYPE505_REG:
                rdata_tmp = jump_type505_reg;
            JUMP_TYPE506_REG:
                rdata_tmp = jump_type506_reg;
            JUMP_TYPE507_REG:
                rdata_tmp = jump_type507_reg;
            JUMP_TYPE508_REG:
                rdata_tmp = jump_type508_reg;
            JUMP_TYPE509_REG:
                rdata_tmp = jump_type509_reg;
            JUMP_TYPE510_REG:
                rdata_tmp = jump_type510_reg;
            JUMP_TYPE511_REG:
                rdata_tmp = jump_type511_reg;
            default:
                rdata_tmp = 32'h0;
        endcase
    end
    else
        rdata_tmp = 32'h0;
end

always @ ( posedge clk or negedge rst_n)
begin
    if( ~rst_n )
        rdata <= 32'h0;
    else if ( ren )
        rdata <= rdata_tmp;
end


endmodule
