//////////////////////////////////////////////////////////////////////////////////
// Description:
//////////////////////////////////////////////////////////////////////////////////

module pdec_rom_stage
#(parameter D=16384,
  parameter W=32,
  parameter RD_TYPE=0) //0=delay address by 1T;1=delay rdata
(
  input                 clk,
  input                 ce,   //high active
  input                 we,   //high active
  input  [$clog2(D)-1:0]addr,
  input  [W-1:0]        wdata,
  output [W-1:0]        rdata
);

  wire [W-1:0] mem[0:D-1]/*synthesis syn_ramstyle="block_ram" */;
  //----intial
  assign mem[0   ] = 5'h18 ; 
  assign mem[1   ] = 5'h17 ;
  assign mem[2   ] = 5'h16 ;
  assign mem[3   ] = 5'h15 ;
  assign mem[4   ] = 5'h14 ;
  assign mem[5   ] = 5'h13 ;
  assign mem[6   ] = 5'h12 ;
  assign mem[7   ] = 5'h11 ;
  assign mem[8   ] = 5'h10 ;
  assign mem[9   ] = 5'h00 ;
  assign mem[10  ] = 5'h01 ;
  assign mem[11  ] = 5'h10 ;
  assign mem[12  ] = 5'h00 ;
  assign mem[13  ] = 5'h02 ;
  assign mem[14  ] = 5'h11 ;
  assign mem[15  ] = 5'h10 ;
  assign mem[16  ] = 5'h00 ;
  assign mem[17  ] = 5'h01 ;
  assign mem[18  ] = 5'h10 ;
  assign mem[19  ] = 5'h00 ;
  assign mem[20  ] = 5'h03 ;
  assign mem[21  ] = 5'h12 ;
  assign mem[22  ] = 5'h11 ;
  assign mem[23  ] = 5'h10 ;
  assign mem[24  ] = 5'h00 ;
  assign mem[25  ] = 5'h01 ;
  assign mem[26  ] = 5'h10 ;
  assign mem[27  ] = 5'h00 ;
  assign mem[28  ] = 5'h02 ;
  assign mem[29  ] = 5'h11 ;
  assign mem[30  ] = 5'h10 ;
  assign mem[31  ] = 5'h00 ;
  assign mem[32  ] = 5'h01 ;
  assign mem[33  ] = 5'h10 ;
  assign mem[34  ] = 5'h00 ;
  assign mem[35  ] = 5'h04 ;
  assign mem[36  ] = 5'h13 ;
  assign mem[37  ] = 5'h12 ;
  assign mem[38  ] = 5'h11 ;
  assign mem[39  ] = 5'h10 ;
  assign mem[40  ] = 5'h00 ;
  assign mem[41  ] = 5'h01 ;
  assign mem[42  ] = 5'h10 ;
  assign mem[43  ] = 5'h00 ;
  assign mem[44  ] = 5'h02 ;
  assign mem[45  ] = 5'h11 ;
  assign mem[46  ] = 5'h10 ;
  assign mem[47  ] = 5'h00 ;
  assign mem[48  ] = 5'h01 ;
  assign mem[49  ] = 5'h10 ;
  assign mem[50  ] = 5'h00 ;
  assign mem[51  ] = 5'h03 ;
  assign mem[52  ] = 5'h12 ;
  assign mem[53  ] = 5'h11 ;
  assign mem[54  ] = 5'h10 ;
  assign mem[55  ] = 5'h00 ;
  assign mem[56  ] = 5'h01 ;
  assign mem[57  ] = 5'h10 ;
  assign mem[58  ] = 5'h00 ;
  assign mem[59  ] = 5'h02 ;
  assign mem[60  ] = 5'h11 ;
  assign mem[61  ] = 5'h10 ;
  assign mem[62  ] = 5'h00 ;
  assign mem[63  ] = 5'h01 ;
  assign mem[64  ] = 5'h10 ;
  assign mem[65  ] = 5'h00 ;
  assign mem[66  ] = 5'h05 ;
  assign mem[67  ] = 5'h14 ;
  assign mem[68  ] = 5'h13 ;
  assign mem[69  ] = 5'h12 ;
  assign mem[70  ] = 5'h11 ;
  assign mem[71  ] = 5'h10 ;
  assign mem[72  ] = 5'h00 ;
  assign mem[73  ] = 5'h01 ;
  assign mem[74  ] = 5'h10 ;
  assign mem[75  ] = 5'h00 ;
  assign mem[76  ] = 5'h02 ;
  assign mem[77  ] = 5'h11 ;
  assign mem[78  ] = 5'h10 ;
  assign mem[79  ] = 5'h00 ;
  assign mem[80  ] = 5'h01 ;
  assign mem[81  ] = 5'h10 ;
  assign mem[82  ] = 5'h00 ;
  assign mem[83  ] = 5'h03 ;
  assign mem[84  ] = 5'h12 ;
  assign mem[85  ] = 5'h11 ;
  assign mem[86  ] = 5'h10 ;
  assign mem[87  ] = 5'h00 ;
  assign mem[88  ] = 5'h01 ;
  assign mem[89  ] = 5'h10 ;
  assign mem[90  ] = 5'h00 ;
  assign mem[91  ] = 5'h02 ;
  assign mem[92  ] = 5'h11 ;
  assign mem[93  ] = 5'h10 ;
  assign mem[94  ] = 5'h00 ;
  assign mem[95  ] = 5'h01 ;
  assign mem[96  ] = 5'h10 ;
  assign mem[97  ] = 5'h00 ;
  assign mem[98  ] = 5'h04 ;
  assign mem[99  ] = 5'h13 ;
  assign mem[100 ] = 5'h12 ;
  assign mem[101 ] = 5'h11 ;
  assign mem[102 ] = 5'h10 ;
  assign mem[103 ] = 5'h00 ;
  assign mem[104 ] = 5'h01 ;
  assign mem[105 ] = 5'h10 ;
  assign mem[106 ] = 5'h00 ;
  assign mem[107 ] = 5'h02 ;
  assign mem[108 ] = 5'h11 ;
  assign mem[109 ] = 5'h10 ;
  assign mem[110 ] = 5'h00 ;
  assign mem[111 ] = 5'h01 ;
  assign mem[112 ] = 5'h10 ;
  assign mem[113 ] = 5'h00 ;
  assign mem[114 ] = 5'h03 ;
  assign mem[115 ] = 5'h12 ;
  assign mem[116 ] = 5'h11 ;
  assign mem[117 ] = 5'h10 ;
  assign mem[118 ] = 5'h00 ;
  assign mem[119 ] = 5'h01 ;
  assign mem[120 ] = 5'h10 ;
  assign mem[121 ] = 5'h00 ;
  assign mem[122 ] = 5'h02 ;
  assign mem[123 ] = 5'h11 ;
  assign mem[124 ] = 5'h10 ;
  assign mem[125 ] = 5'h00 ;
  assign mem[126 ] = 5'h01 ;
  assign mem[127 ] = 5'h10 ;
  assign mem[128 ] = 5'h00 ;
  assign mem[129 ] = 5'h06 ;
  assign mem[130 ] = 5'h15 ;
  assign mem[131 ] = 5'h14 ;
  assign mem[132 ] = 5'h13 ;
  assign mem[133 ] = 5'h12 ;
  assign mem[134 ] = 5'h11 ;
  assign mem[135 ] = 5'h10 ;
  assign mem[136 ] = 5'h00 ;
  assign mem[137 ] = 5'h01 ;
  assign mem[138 ] = 5'h10 ;
  assign mem[139 ] = 5'h00 ;
  assign mem[140 ] = 5'h02 ;
  assign mem[141 ] = 5'h11 ;
  assign mem[142 ] = 5'h10 ;
  assign mem[143 ] = 5'h00 ;
  assign mem[144 ] = 5'h01 ;
  assign mem[145 ] = 5'h10 ;
  assign mem[146 ] = 5'h00 ;
  assign mem[147 ] = 5'h03 ;
  assign mem[148 ] = 5'h12 ;
  assign mem[149 ] = 5'h11 ;
  assign mem[150 ] = 5'h10 ;
  assign mem[151 ] = 5'h00 ;
  assign mem[152 ] = 5'h01 ;
  assign mem[153 ] = 5'h10 ;
  assign mem[154 ] = 5'h00 ;
  assign mem[155 ] = 5'h02 ;
  assign mem[156 ] = 5'h11 ;
  assign mem[157 ] = 5'h10 ;
  assign mem[158 ] = 5'h00 ;
  assign mem[159 ] = 5'h01 ;
  assign mem[160 ] = 5'h10 ;
  assign mem[161 ] = 5'h00 ;
  assign mem[162 ] = 5'h04 ;
  assign mem[163 ] = 5'h13 ;
  assign mem[164 ] = 5'h12 ;
  assign mem[165 ] = 5'h11 ;
  assign mem[166 ] = 5'h10 ;
  assign mem[167 ] = 5'h00 ;
  assign mem[168 ] = 5'h01 ;
  assign mem[169 ] = 5'h10 ;
  assign mem[170 ] = 5'h00 ;
  assign mem[171 ] = 5'h02 ;
  assign mem[172 ] = 5'h11 ;
  assign mem[173 ] = 5'h10 ;
  assign mem[174 ] = 5'h00 ;
  assign mem[175 ] = 5'h01 ;
  assign mem[176 ] = 5'h10 ;
  assign mem[177 ] = 5'h00 ;
  assign mem[178 ] = 5'h03 ;
  assign mem[179 ] = 5'h12 ;
  assign mem[180 ] = 5'h11 ;
  assign mem[181 ] = 5'h10 ;
  assign mem[182 ] = 5'h00 ;
  assign mem[183 ] = 5'h01 ;
  assign mem[184 ] = 5'h10 ;
  assign mem[185 ] = 5'h00 ;
  assign mem[186 ] = 5'h02 ;
  assign mem[187 ] = 5'h11 ;
  assign mem[188 ] = 5'h10 ;
  assign mem[189 ] = 5'h00 ;
  assign mem[190 ] = 5'h01 ;
  assign mem[191 ] = 5'h10 ;
  assign mem[192 ] = 5'h00 ;
  assign mem[193 ] = 5'h05 ;
  assign mem[194 ] = 5'h14 ;
  assign mem[195 ] = 5'h13 ;
  assign mem[196 ] = 5'h12 ;
  assign mem[197 ] = 5'h11 ;
  assign mem[198 ] = 5'h10 ;
  assign mem[199 ] = 5'h00 ;
  assign mem[200 ] = 5'h01 ;
  assign mem[201 ] = 5'h10 ;
  assign mem[202 ] = 5'h00 ;
  assign mem[203 ] = 5'h02 ;
  assign mem[204 ] = 5'h11 ;
  assign mem[205 ] = 5'h10 ;
  assign mem[206 ] = 5'h00 ;
  assign mem[207 ] = 5'h01 ;
  assign mem[208 ] = 5'h10 ;
  assign mem[209 ] = 5'h00 ;
  assign mem[210 ] = 5'h03 ;
  assign mem[211 ] = 5'h12 ;
  assign mem[212 ] = 5'h11 ;
  assign mem[213 ] = 5'h10 ;
  assign mem[214 ] = 5'h00 ;
  assign mem[215 ] = 5'h01 ;
  assign mem[216 ] = 5'h10 ;
  assign mem[217 ] = 5'h00 ;
  assign mem[218 ] = 5'h02 ;
  assign mem[219 ] = 5'h11 ;
  assign mem[220 ] = 5'h10 ;
  assign mem[221 ] = 5'h00 ;
  assign mem[222 ] = 5'h01 ;
  assign mem[223 ] = 5'h10 ;
  assign mem[224 ] = 5'h00 ;
  assign mem[225 ] = 5'h04 ;
  assign mem[226 ] = 5'h13 ;
  assign mem[227 ] = 5'h12 ;
  assign mem[228 ] = 5'h11 ;
  assign mem[229 ] = 5'h10 ;
  assign mem[230 ] = 5'h00 ;
  assign mem[231 ] = 5'h01 ;
  assign mem[232 ] = 5'h10 ;
  assign mem[233 ] = 5'h00 ;
  assign mem[234 ] = 5'h02 ;
  assign mem[235 ] = 5'h11 ;
  assign mem[236 ] = 5'h10 ;
  assign mem[237 ] = 5'h00 ;
  assign mem[238 ] = 5'h01 ;
  assign mem[239 ] = 5'h10 ;
  assign mem[240 ] = 5'h00 ;
  assign mem[241 ] = 5'h03 ;
  assign mem[242 ] = 5'h12 ;
  assign mem[243 ] = 5'h11 ;
  assign mem[244 ] = 5'h10 ;
  assign mem[245 ] = 5'h00 ;
  assign mem[246 ] = 5'h01 ;
  assign mem[247 ] = 5'h10 ;
  assign mem[248 ] = 5'h00 ;
  assign mem[249 ] = 5'h02 ;
  assign mem[250 ] = 5'h11 ;
  assign mem[251 ] = 5'h10 ;
  assign mem[252 ] = 5'h00 ;
  assign mem[253 ] = 5'h01 ;
  assign mem[254 ] = 5'h10 ;
  assign mem[255 ] = 5'h00 ;
  assign mem[256 ] = 5'h07 ;
  assign mem[257 ] = 5'h16 ;
  assign mem[258 ] = 5'h15 ;
  assign mem[259 ] = 5'h14 ;
  assign mem[260 ] = 5'h13 ;
  assign mem[261 ] = 5'h12 ;
  assign mem[262 ] = 5'h11 ;
  assign mem[263 ] = 5'h10 ;
  assign mem[264 ] = 5'h00 ;
  assign mem[265 ] = 5'h01 ;
  assign mem[266 ] = 5'h10 ;
  assign mem[267 ] = 5'h00 ;
  assign mem[268 ] = 5'h02 ;
  assign mem[269 ] = 5'h11 ;
  assign mem[270 ] = 5'h10 ;
  assign mem[271 ] = 5'h00 ;
  assign mem[272 ] = 5'h01 ;
  assign mem[273 ] = 5'h10 ;
  assign mem[274 ] = 5'h00 ;
  assign mem[275 ] = 5'h03 ;
  assign mem[276 ] = 5'h12 ;
  assign mem[277 ] = 5'h11 ;
  assign mem[278 ] = 5'h10 ;
  assign mem[279 ] = 5'h00 ;
  assign mem[280 ] = 5'h01 ;
  assign mem[281 ] = 5'h10 ;
  assign mem[282 ] = 5'h00 ;
  assign mem[283 ] = 5'h02 ;
  assign mem[284 ] = 5'h11 ;
  assign mem[285 ] = 5'h10 ;
  assign mem[286 ] = 5'h00 ;
  assign mem[287 ] = 5'h01 ;
  assign mem[288 ] = 5'h10 ;
  assign mem[289 ] = 5'h00 ;
  assign mem[290 ] = 5'h04 ;
  assign mem[291 ] = 5'h13 ;
  assign mem[292 ] = 5'h12 ;
  assign mem[293 ] = 5'h11 ;
  assign mem[294 ] = 5'h10 ;
  assign mem[295 ] = 5'h00 ;
  assign mem[296 ] = 5'h01 ;
  assign mem[297 ] = 5'h10 ;
  assign mem[298 ] = 5'h00 ;
  assign mem[299 ] = 5'h02 ;
  assign mem[300 ] = 5'h11 ;
  assign mem[301 ] = 5'h10 ;
  assign mem[302 ] = 5'h00 ;
  assign mem[303 ] = 5'h01 ;
  assign mem[304 ] = 5'h10 ;
  assign mem[305 ] = 5'h00 ;
  assign mem[306 ] = 5'h03 ;
  assign mem[307 ] = 5'h12 ;
  assign mem[308 ] = 5'h11 ;
  assign mem[309 ] = 5'h10 ;
  assign mem[310 ] = 5'h00 ;
  assign mem[311 ] = 5'h01 ;
  assign mem[312 ] = 5'h10 ;
  assign mem[313 ] = 5'h00 ;
  assign mem[314 ] = 5'h02 ;
  assign mem[315 ] = 5'h11 ;
  assign mem[316 ] = 5'h10 ;
  assign mem[317 ] = 5'h00 ;
  assign mem[318 ] = 5'h01 ;
  assign mem[319 ] = 5'h10 ;
  assign mem[320 ] = 5'h00 ;
  assign mem[321 ] = 5'h05 ;
  assign mem[322 ] = 5'h14 ;
  assign mem[323 ] = 5'h13 ;
  assign mem[324 ] = 5'h12 ;
  assign mem[325 ] = 5'h11 ;
  assign mem[326 ] = 5'h10 ;
  assign mem[327 ] = 5'h00 ;
  assign mem[328 ] = 5'h01 ;
  assign mem[329 ] = 5'h10 ;
  assign mem[330 ] = 5'h00 ;
  assign mem[331 ] = 5'h02 ;
  assign mem[332 ] = 5'h11 ;
  assign mem[333 ] = 5'h10 ;
  assign mem[334 ] = 5'h00 ;
  assign mem[335 ] = 5'h01 ;
  assign mem[336 ] = 5'h10 ;
  assign mem[337 ] = 5'h00 ;
  assign mem[338 ] = 5'h03 ;
  assign mem[339 ] = 5'h12 ;
  assign mem[340 ] = 5'h11 ;
  assign mem[341 ] = 5'h10 ;
  assign mem[342 ] = 5'h00 ;
  assign mem[343 ] = 5'h01 ;
  assign mem[344 ] = 5'h10 ;
  assign mem[345 ] = 5'h00 ;
  assign mem[346 ] = 5'h02 ;
  assign mem[347 ] = 5'h11 ;
  assign mem[348 ] = 5'h10 ;
  assign mem[349 ] = 5'h00 ;
  assign mem[350 ] = 5'h01 ;
  assign mem[351 ] = 5'h10 ;
  assign mem[352 ] = 5'h00 ;
  assign mem[353 ] = 5'h04 ;
  assign mem[354 ] = 5'h13 ;
  assign mem[355 ] = 5'h12 ;
  assign mem[356 ] = 5'h11 ;
  assign mem[357 ] = 5'h10 ;
  assign mem[358 ] = 5'h00 ;
  assign mem[359 ] = 5'h01 ;
  assign mem[360 ] = 5'h10 ;
  assign mem[361 ] = 5'h00 ;
  assign mem[362 ] = 5'h02 ;
  assign mem[363 ] = 5'h11 ;
  assign mem[364 ] = 5'h10 ;
  assign mem[365 ] = 5'h00 ;
  assign mem[366 ] = 5'h01 ;
  assign mem[367 ] = 5'h10 ;
  assign mem[368 ] = 5'h00 ;
  assign mem[369 ] = 5'h03 ;
  assign mem[370 ] = 5'h12 ;
  assign mem[371 ] = 5'h11 ;
  assign mem[372 ] = 5'h10 ;
  assign mem[373 ] = 5'h00 ;
  assign mem[374 ] = 5'h01 ;
  assign mem[375 ] = 5'h10 ;
  assign mem[376 ] = 5'h00 ;
  assign mem[377 ] = 5'h02 ;
  assign mem[378 ] = 5'h11 ;
  assign mem[379 ] = 5'h10 ;
  assign mem[380 ] = 5'h00 ;
  assign mem[381 ] = 5'h01 ;
  assign mem[382 ] = 5'h10 ;
  assign mem[383 ] = 5'h00 ;
  assign mem[384 ] = 5'h06 ;
  assign mem[385 ] = 5'h15 ;
  assign mem[386 ] = 5'h14 ;
  assign mem[387 ] = 5'h13 ;
  assign mem[388 ] = 5'h12 ;
  assign mem[389 ] = 5'h11 ;
  assign mem[390 ] = 5'h10 ;
  assign mem[391 ] = 5'h00 ;
  assign mem[392 ] = 5'h01 ;
  assign mem[393 ] = 5'h10 ;
  assign mem[394 ] = 5'h00 ;
  assign mem[395 ] = 5'h02 ;
  assign mem[396 ] = 5'h11 ;
  assign mem[397 ] = 5'h10 ;
  assign mem[398 ] = 5'h00 ;
  assign mem[399 ] = 5'h01 ;
  assign mem[400 ] = 5'h10 ;
  assign mem[401 ] = 5'h00 ;
  assign mem[402 ] = 5'h03 ;
  assign mem[403 ] = 5'h12 ;
  assign mem[404 ] = 5'h11 ;
  assign mem[405 ] = 5'h10 ;
  assign mem[406 ] = 5'h00 ;
  assign mem[407 ] = 5'h01 ;
  assign mem[408 ] = 5'h10 ;
  assign mem[409 ] = 5'h00 ;
  assign mem[410 ] = 5'h02 ;
  assign mem[411 ] = 5'h11 ;
  assign mem[412 ] = 5'h10 ;
  assign mem[413 ] = 5'h00 ;
  assign mem[414 ] = 5'h01 ;
  assign mem[415 ] = 5'h10 ;
  assign mem[416 ] = 5'h00 ;
  assign mem[417 ] = 5'h04 ;
  assign mem[418 ] = 5'h13 ;
  assign mem[419 ] = 5'h12 ;
  assign mem[420 ] = 5'h11 ;
  assign mem[421 ] = 5'h10 ;
  assign mem[422 ] = 5'h00 ;
  assign mem[423 ] = 5'h01 ;
  assign mem[424 ] = 5'h10 ;
  assign mem[425 ] = 5'h00 ;
  assign mem[426 ] = 5'h02 ;
  assign mem[427 ] = 5'h11 ;
  assign mem[428 ] = 5'h10 ;
  assign mem[429 ] = 5'h00 ;
  assign mem[430 ] = 5'h01 ;
  assign mem[431 ] = 5'h10 ;
  assign mem[432 ] = 5'h00 ;
  assign mem[433 ] = 5'h03 ;
  assign mem[434 ] = 5'h12 ;
  assign mem[435 ] = 5'h11 ;
  assign mem[436 ] = 5'h10 ;
  assign mem[437 ] = 5'h00 ;
  assign mem[438 ] = 5'h01 ;
  assign mem[439 ] = 5'h10 ;
  assign mem[440 ] = 5'h00 ;
  assign mem[441 ] = 5'h02 ;
  assign mem[442 ] = 5'h11 ;
  assign mem[443 ] = 5'h10 ;
  assign mem[444 ] = 5'h00 ;
  assign mem[445 ] = 5'h01 ;
  assign mem[446 ] = 5'h10 ;
  assign mem[447 ] = 5'h00 ;
  assign mem[448 ] = 5'h05 ;
  assign mem[449 ] = 5'h14 ;
  assign mem[450 ] = 5'h13 ;
  assign mem[451 ] = 5'h12 ;
  assign mem[452 ] = 5'h11 ;
  assign mem[453 ] = 5'h10 ;
  assign mem[454 ] = 5'h00 ;
  assign mem[455 ] = 5'h01 ;
  assign mem[456 ] = 5'h10 ;
  assign mem[457 ] = 5'h00 ;
  assign mem[458 ] = 5'h02 ;
  assign mem[459 ] = 5'h11 ;
  assign mem[460 ] = 5'h10 ;
  assign mem[461 ] = 5'h00 ;
  assign mem[462 ] = 5'h01 ;
  assign mem[463 ] = 5'h10 ;
  assign mem[464 ] = 5'h00 ;
  assign mem[465 ] = 5'h03 ;
  assign mem[466 ] = 5'h12 ;
  assign mem[467 ] = 5'h11 ;
  assign mem[468 ] = 5'h10 ;
  assign mem[469 ] = 5'h00 ;
  assign mem[470 ] = 5'h01 ;
  assign mem[471 ] = 5'h10 ;
  assign mem[472 ] = 5'h00 ;
  assign mem[473 ] = 5'h02 ;
  assign mem[474 ] = 5'h11 ;
  assign mem[475 ] = 5'h10 ;
  assign mem[476 ] = 5'h00 ;
  assign mem[477 ] = 5'h01 ;
  assign mem[478 ] = 5'h10 ;
  assign mem[479 ] = 5'h00 ;
  assign mem[480 ] = 5'h04 ;
  assign mem[481 ] = 5'h13 ;
  assign mem[482 ] = 5'h12 ;
  assign mem[483 ] = 5'h11 ;
  assign mem[484 ] = 5'h10 ;
  assign mem[485 ] = 5'h00 ;
  assign mem[486 ] = 5'h01 ;
  assign mem[487 ] = 5'h10 ;
  assign mem[488 ] = 5'h00 ;
  assign mem[489 ] = 5'h02 ;
  assign mem[490 ] = 5'h11 ;
  assign mem[491 ] = 5'h10 ;
  assign mem[492 ] = 5'h00 ;
  assign mem[493 ] = 5'h01 ;
  assign mem[494 ] = 5'h10 ;
  assign mem[495 ] = 5'h00 ;
  assign mem[496 ] = 5'h03 ;
  assign mem[497 ] = 5'h12 ;
  assign mem[498 ] = 5'h11 ;
  assign mem[499 ] = 5'h10 ;
  assign mem[500 ] = 5'h00 ;
  assign mem[501 ] = 5'h01 ;
  assign mem[502 ] = 5'h10 ;
  assign mem[503 ] = 5'h00 ;
  assign mem[504 ] = 5'h02 ;
  assign mem[505 ] = 5'h11 ;
  assign mem[506 ] = 5'h10 ;
  assign mem[507 ] = 5'h00 ;
  assign mem[508 ] = 5'h01 ;
  assign mem[509 ] = 5'h10 ;
  assign mem[510 ] = 5'h00 ;
  assign mem[511 ] = 5'h08 ;
  assign mem[512 ] = 5'h17 ;
  assign mem[513 ] = 5'h16 ;
  assign mem[514 ] = 5'h15 ;
  assign mem[515 ] = 5'h14 ;
  assign mem[516 ] = 5'h13 ;
  assign mem[517 ] = 5'h12 ;
  assign mem[518 ] = 5'h11 ;
  assign mem[519 ] = 5'h10 ;
  assign mem[520 ] = 5'h00 ;
  assign mem[521 ] = 5'h01 ;
  assign mem[522 ] = 5'h10 ;
  assign mem[523 ] = 5'h00 ;
  assign mem[524 ] = 5'h02 ;
  assign mem[525 ] = 5'h11 ;
  assign mem[526 ] = 5'h10 ;
  assign mem[527 ] = 5'h00 ;
  assign mem[528 ] = 5'h01 ;
  assign mem[529 ] = 5'h10 ;
  assign mem[530 ] = 5'h00 ;
  assign mem[531 ] = 5'h03 ;
  assign mem[532 ] = 5'h12 ;
  assign mem[533 ] = 5'h11 ;
  assign mem[534 ] = 5'h10 ;
  assign mem[535 ] = 5'h00 ;
  assign mem[536 ] = 5'h01 ;
  assign mem[537 ] = 5'h10 ;
  assign mem[538 ] = 5'h00 ;
  assign mem[539 ] = 5'h02 ;
  assign mem[540 ] = 5'h11 ;
  assign mem[541 ] = 5'h10 ;
  assign mem[542 ] = 5'h00 ;
  assign mem[543 ] = 5'h01 ;
  assign mem[544 ] = 5'h10 ;
  assign mem[545 ] = 5'h00 ;
  assign mem[546 ] = 5'h04 ;
  assign mem[547 ] = 5'h13 ;
  assign mem[548 ] = 5'h12 ;
  assign mem[549 ] = 5'h11 ;
  assign mem[550 ] = 5'h10 ;
  assign mem[551 ] = 5'h00 ;
  assign mem[552 ] = 5'h01 ;
  assign mem[553 ] = 5'h10 ;
  assign mem[554 ] = 5'h00 ;
  assign mem[555 ] = 5'h02 ;
  assign mem[556 ] = 5'h11 ;
  assign mem[557 ] = 5'h10 ;
  assign mem[558 ] = 5'h00 ;
  assign mem[559 ] = 5'h01 ;
  assign mem[560 ] = 5'h10 ;
  assign mem[561 ] = 5'h00 ;
  assign mem[562 ] = 5'h03 ;
  assign mem[563 ] = 5'h12 ;
  assign mem[564 ] = 5'h11 ;
  assign mem[565 ] = 5'h10 ;
  assign mem[566 ] = 5'h00 ;
  assign mem[567 ] = 5'h01 ;
  assign mem[568 ] = 5'h10 ;
  assign mem[569 ] = 5'h00 ;
  assign mem[570 ] = 5'h02 ;
  assign mem[571 ] = 5'h11 ;
  assign mem[572 ] = 5'h10 ;
  assign mem[573 ] = 5'h00 ;
  assign mem[574 ] = 5'h01 ;
  assign mem[575 ] = 5'h10 ;
  assign mem[576 ] = 5'h00 ;
  assign mem[577 ] = 5'h05 ;
  assign mem[578 ] = 5'h14 ;
  assign mem[579 ] = 5'h13 ;
  assign mem[580 ] = 5'h12 ;
  assign mem[581 ] = 5'h11 ;
  assign mem[582 ] = 5'h10 ;
  assign mem[583 ] = 5'h00 ;
  assign mem[584 ] = 5'h01 ;
  assign mem[585 ] = 5'h10 ;
  assign mem[586 ] = 5'h00 ;
  assign mem[587 ] = 5'h02 ;
  assign mem[588 ] = 5'h11 ;
  assign mem[589 ] = 5'h10 ;
  assign mem[590 ] = 5'h00 ;
  assign mem[591 ] = 5'h01 ;
  assign mem[592 ] = 5'h10 ;
  assign mem[593 ] = 5'h00 ;
  assign mem[594 ] = 5'h03 ;
  assign mem[595 ] = 5'h12 ;
  assign mem[596 ] = 5'h11 ;
  assign mem[597 ] = 5'h10 ;
  assign mem[598 ] = 5'h00 ;
  assign mem[599 ] = 5'h01 ;
  assign mem[600 ] = 5'h10 ;
  assign mem[601 ] = 5'h00 ;
  assign mem[602 ] = 5'h02 ;
  assign mem[603 ] = 5'h11 ;
  assign mem[604 ] = 5'h10 ;
  assign mem[605 ] = 5'h00 ;
  assign mem[606 ] = 5'h01 ;
  assign mem[607 ] = 5'h10 ;
  assign mem[608 ] = 5'h00 ;
  assign mem[609 ] = 5'h04 ;
  assign mem[610 ] = 5'h13 ;
  assign mem[611 ] = 5'h12 ;
  assign mem[612 ] = 5'h11 ;
  assign mem[613 ] = 5'h10 ;
  assign mem[614 ] = 5'h00 ;
  assign mem[615 ] = 5'h01 ;
  assign mem[616 ] = 5'h10 ;
  assign mem[617 ] = 5'h00 ;
  assign mem[618 ] = 5'h02 ;
  assign mem[619 ] = 5'h11 ;
  assign mem[620 ] = 5'h10 ;
  assign mem[621 ] = 5'h00 ;
  assign mem[622 ] = 5'h01 ;
  assign mem[623 ] = 5'h10 ;
  assign mem[624 ] = 5'h00 ;
  assign mem[625 ] = 5'h03 ;
  assign mem[626 ] = 5'h12 ;
  assign mem[627 ] = 5'h11 ;
  assign mem[628 ] = 5'h10 ;
  assign mem[629 ] = 5'h00 ;
  assign mem[630 ] = 5'h01 ;
  assign mem[631 ] = 5'h10 ;
  assign mem[632 ] = 5'h00 ;
  assign mem[633 ] = 5'h02 ;
  assign mem[634 ] = 5'h11 ;
  assign mem[635 ] = 5'h10 ;
  assign mem[636 ] = 5'h00 ;
  assign mem[637 ] = 5'h01 ;
  assign mem[638 ] = 5'h10 ;
  assign mem[639 ] = 5'h00 ;
  assign mem[640 ] = 5'h06 ;
  assign mem[641 ] = 5'h15 ;
  assign mem[642 ] = 5'h14 ;
  assign mem[643 ] = 5'h13 ;
  assign mem[644 ] = 5'h12 ;
  assign mem[645 ] = 5'h11 ;
  assign mem[646 ] = 5'h10 ;
  assign mem[647 ] = 5'h00 ;
  assign mem[648 ] = 5'h01 ;
  assign mem[649 ] = 5'h10 ;
  assign mem[650 ] = 5'h00 ;
  assign mem[651 ] = 5'h02 ;
  assign mem[652 ] = 5'h11 ;
  assign mem[653 ] = 5'h10 ;
  assign mem[654 ] = 5'h00 ;
  assign mem[655 ] = 5'h01 ;
  assign mem[656 ] = 5'h10 ;
  assign mem[657 ] = 5'h00 ;
  assign mem[658 ] = 5'h03 ;
  assign mem[659 ] = 5'h12 ;
  assign mem[660 ] = 5'h11 ;
  assign mem[661 ] = 5'h10 ;
  assign mem[662 ] = 5'h00 ;
  assign mem[663 ] = 5'h01 ;
  assign mem[664 ] = 5'h10 ;
  assign mem[665 ] = 5'h00 ;
  assign mem[666 ] = 5'h02 ;
  assign mem[667 ] = 5'h11 ;
  assign mem[668 ] = 5'h10 ;
  assign mem[669 ] = 5'h00 ;
  assign mem[670 ] = 5'h01 ;
  assign mem[671 ] = 5'h10 ;
  assign mem[672 ] = 5'h00 ;
  assign mem[673 ] = 5'h04 ;
  assign mem[674 ] = 5'h13 ;
  assign mem[675 ] = 5'h12 ;
  assign mem[676 ] = 5'h11 ;
  assign mem[677 ] = 5'h10 ;
  assign mem[678 ] = 5'h00 ;
  assign mem[679 ] = 5'h01 ;
  assign mem[680 ] = 5'h10 ;
  assign mem[681 ] = 5'h00 ;
  assign mem[682 ] = 5'h02 ;
  assign mem[683 ] = 5'h11 ;
  assign mem[684 ] = 5'h10 ;
  assign mem[685 ] = 5'h00 ;
  assign mem[686 ] = 5'h01 ;
  assign mem[687 ] = 5'h10 ;
  assign mem[688 ] = 5'h00 ;
  assign mem[689 ] = 5'h03 ;
  assign mem[690 ] = 5'h12 ;
  assign mem[691 ] = 5'h11 ;
  assign mem[692 ] = 5'h10 ;
  assign mem[693 ] = 5'h00 ;
  assign mem[694 ] = 5'h01 ;
  assign mem[695 ] = 5'h10 ;
  assign mem[696 ] = 5'h00 ;
  assign mem[697 ] = 5'h02 ;
  assign mem[698 ] = 5'h11 ;
  assign mem[699 ] = 5'h10 ;
  assign mem[700 ] = 5'h00 ;
  assign mem[701 ] = 5'h01 ;
  assign mem[702 ] = 5'h10 ;
  assign mem[703 ] = 5'h00 ;
  assign mem[704 ] = 5'h05 ;
  assign mem[705 ] = 5'h14 ;
  assign mem[706 ] = 5'h13 ;
  assign mem[707 ] = 5'h12 ;
  assign mem[708 ] = 5'h11 ;
  assign mem[709 ] = 5'h10 ;
  assign mem[710 ] = 5'h00 ;
  assign mem[711 ] = 5'h01 ;
  assign mem[712 ] = 5'h10 ;
  assign mem[713 ] = 5'h00 ;
  assign mem[714 ] = 5'h02 ;
  assign mem[715 ] = 5'h11 ;
  assign mem[716 ] = 5'h10 ;
  assign mem[717 ] = 5'h00 ;
  assign mem[718 ] = 5'h01 ;
  assign mem[719 ] = 5'h10 ;
  assign mem[720 ] = 5'h00 ;
  assign mem[721 ] = 5'h03 ;
  assign mem[722 ] = 5'h12 ;
  assign mem[723 ] = 5'h11 ;
  assign mem[724 ] = 5'h10 ;
  assign mem[725 ] = 5'h00 ;
  assign mem[726 ] = 5'h01 ;
  assign mem[727 ] = 5'h10 ;
  assign mem[728 ] = 5'h00 ;
  assign mem[729 ] = 5'h02 ;
  assign mem[730 ] = 5'h11 ;
  assign mem[731 ] = 5'h10 ;
  assign mem[732 ] = 5'h00 ;
  assign mem[733 ] = 5'h01 ;
  assign mem[734 ] = 5'h10 ;
  assign mem[735 ] = 5'h00 ;
  assign mem[736 ] = 5'h04 ;
  assign mem[737 ] = 5'h13 ;
  assign mem[738 ] = 5'h12 ;
  assign mem[739 ] = 5'h11 ;
  assign mem[740 ] = 5'h10 ;
  assign mem[741 ] = 5'h00 ;
  assign mem[742 ] = 5'h01 ;
  assign mem[743 ] = 5'h10 ;
  assign mem[744 ] = 5'h00 ;
  assign mem[745 ] = 5'h02 ;
  assign mem[746 ] = 5'h11 ;
  assign mem[747 ] = 5'h10 ;
  assign mem[748 ] = 5'h00 ;
  assign mem[749 ] = 5'h01 ;
  assign mem[750 ] = 5'h10 ;
  assign mem[751 ] = 5'h00 ;
  assign mem[752 ] = 5'h03 ;
  assign mem[753 ] = 5'h12 ;
  assign mem[754 ] = 5'h11 ;
  assign mem[755 ] = 5'h10 ;
  assign mem[756 ] = 5'h00 ;
  assign mem[757 ] = 5'h01 ;
  assign mem[758 ] = 5'h10 ;
  assign mem[759 ] = 5'h00 ;
  assign mem[760 ] = 5'h02 ;
  assign mem[761 ] = 5'h11 ;
  assign mem[762 ] = 5'h10 ;
  assign mem[763 ] = 5'h00 ;
  assign mem[764 ] = 5'h01 ;
  assign mem[765 ] = 5'h10 ;
  assign mem[766 ] = 5'h00 ;
  assign mem[767 ] = 5'h07 ;
  assign mem[768 ] = 5'h16 ;
  assign mem[769 ] = 5'h15 ;
  assign mem[770 ] = 5'h14 ;
  assign mem[771 ] = 5'h13 ;
  assign mem[772 ] = 5'h12 ;
  assign mem[773 ] = 5'h11 ;
  assign mem[774 ] = 5'h10 ;
  assign mem[775 ] = 5'h00 ;
  assign mem[776 ] = 5'h01 ;
  assign mem[777 ] = 5'h10 ;
  assign mem[778 ] = 5'h00 ;
  assign mem[779 ] = 5'h02 ;
  assign mem[780 ] = 5'h11 ;
  assign mem[781 ] = 5'h10 ;
  assign mem[782 ] = 5'h00 ;
  assign mem[783 ] = 5'h01 ;
  assign mem[784 ] = 5'h10 ;
  assign mem[785 ] = 5'h00 ;
  assign mem[786 ] = 5'h03 ;
  assign mem[787 ] = 5'h12 ;
  assign mem[788 ] = 5'h11 ;
  assign mem[789 ] = 5'h10 ;
  assign mem[790 ] = 5'h00 ;
  assign mem[791 ] = 5'h01 ;
  assign mem[792 ] = 5'h10 ;
  assign mem[793 ] = 5'h00 ;
  assign mem[794 ] = 5'h02 ;
  assign mem[795 ] = 5'h11 ;
  assign mem[796 ] = 5'h10 ;
  assign mem[797 ] = 5'h00 ;
  assign mem[798 ] = 5'h01 ;
  assign mem[799 ] = 5'h10 ;
  assign mem[800 ] = 5'h00 ;
  assign mem[801 ] = 5'h04 ;
  assign mem[802 ] = 5'h13 ;
  assign mem[803 ] = 5'h12 ;
  assign mem[804 ] = 5'h11 ;
  assign mem[805 ] = 5'h10 ;
  assign mem[806 ] = 5'h00 ;
  assign mem[807 ] = 5'h01 ;
  assign mem[808 ] = 5'h10 ;
  assign mem[809 ] = 5'h00 ;
  assign mem[810 ] = 5'h02 ;
  assign mem[811 ] = 5'h11 ;
  assign mem[812 ] = 5'h10 ;
  assign mem[813 ] = 5'h00 ;
  assign mem[814 ] = 5'h01 ;
  assign mem[815 ] = 5'h10 ;
  assign mem[816 ] = 5'h00 ;
  assign mem[817 ] = 5'h03 ;
  assign mem[818 ] = 5'h12 ;
  assign mem[819 ] = 5'h11 ;
  assign mem[820 ] = 5'h10 ;
  assign mem[821 ] = 5'h00 ;
  assign mem[822 ] = 5'h01 ;
  assign mem[823 ] = 5'h10 ;
  assign mem[824 ] = 5'h00 ;
  assign mem[825 ] = 5'h02 ;
  assign mem[826 ] = 5'h11 ;
  assign mem[827 ] = 5'h10 ;
  assign mem[828 ] = 5'h00 ;
  assign mem[829 ] = 5'h01 ;
  assign mem[830 ] = 5'h10 ;
  assign mem[831 ] = 5'h00 ;
  assign mem[832 ] = 5'h05 ;
  assign mem[833 ] = 5'h14 ;
  assign mem[834 ] = 5'h13 ;
  assign mem[835 ] = 5'h12 ;
  assign mem[836 ] = 5'h11 ;
  assign mem[837 ] = 5'h10 ;
  assign mem[838 ] = 5'h00 ;
  assign mem[839 ] = 5'h01 ;
  assign mem[840 ] = 5'h10 ;
  assign mem[841 ] = 5'h00 ;
  assign mem[842 ] = 5'h02 ;
  assign mem[843 ] = 5'h11 ;
  assign mem[844 ] = 5'h10 ;
  assign mem[845 ] = 5'h00 ;
  assign mem[846 ] = 5'h01 ;
  assign mem[847 ] = 5'h10 ;
  assign mem[848 ] = 5'h00 ;
  assign mem[849 ] = 5'h03 ;
  assign mem[850 ] = 5'h12 ;
  assign mem[851 ] = 5'h11 ;
  assign mem[852 ] = 5'h10 ;
  assign mem[853 ] = 5'h00 ;
  assign mem[854 ] = 5'h01 ;
  assign mem[855 ] = 5'h10 ;
  assign mem[856 ] = 5'h00 ;
  assign mem[857 ] = 5'h02 ;
  assign mem[858 ] = 5'h11 ;
  assign mem[859 ] = 5'h10 ;
  assign mem[860 ] = 5'h00 ;
  assign mem[861 ] = 5'h01 ;
  assign mem[862 ] = 5'h10 ;
  assign mem[863 ] = 5'h00 ;
  assign mem[864 ] = 5'h04 ;
  assign mem[865 ] = 5'h13 ;
  assign mem[866 ] = 5'h12 ;
  assign mem[867 ] = 5'h11 ;
  assign mem[868 ] = 5'h10 ;
  assign mem[869 ] = 5'h00 ;
  assign mem[870 ] = 5'h01 ;
  assign mem[871 ] = 5'h10 ;
  assign mem[872 ] = 5'h00 ;
  assign mem[873 ] = 5'h02 ;
  assign mem[874 ] = 5'h11 ;
  assign mem[875 ] = 5'h10 ;
  assign mem[876 ] = 5'h00 ;
  assign mem[877 ] = 5'h01 ;
  assign mem[878 ] = 5'h10 ;
  assign mem[879 ] = 5'h00 ;
  assign mem[880 ] = 5'h03 ;
  assign mem[881 ] = 5'h12 ;
  assign mem[882 ] = 5'h11 ;
  assign mem[883 ] = 5'h10 ;
  assign mem[884 ] = 5'h00 ;
  assign mem[885 ] = 5'h01 ;
  assign mem[886 ] = 5'h10 ;
  assign mem[887 ] = 5'h00 ;
  assign mem[888 ] = 5'h02 ;
  assign mem[889 ] = 5'h11 ;
  assign mem[890 ] = 5'h10 ;
  assign mem[891 ] = 5'h00 ;
  assign mem[892 ] = 5'h01 ;
  assign mem[893 ] = 5'h10 ;
  assign mem[894 ] = 5'h00 ;
  assign mem[895 ] = 5'h06 ;
  assign mem[896 ] = 5'h15 ;
  assign mem[897 ] = 5'h14 ;
  assign mem[898 ] = 5'h13 ;
  assign mem[899 ] = 5'h12 ;
  assign mem[900 ] = 5'h11 ;
  assign mem[901 ] = 5'h10 ;
  assign mem[902 ] = 5'h00 ;
  assign mem[903 ] = 5'h01 ;
  assign mem[904 ] = 5'h10 ;
  assign mem[905 ] = 5'h00 ;
  assign mem[906 ] = 5'h02 ;
  assign mem[907 ] = 5'h11 ;
  assign mem[908 ] = 5'h10 ;
  assign mem[909 ] = 5'h00 ;
  assign mem[910 ] = 5'h01 ;
  assign mem[911 ] = 5'h10 ;
  assign mem[912 ] = 5'h00 ;
  assign mem[913 ] = 5'h03 ;
  assign mem[914 ] = 5'h12 ;
  assign mem[915 ] = 5'h11 ;
  assign mem[916 ] = 5'h10 ;
  assign mem[917 ] = 5'h00 ;
  assign mem[918 ] = 5'h01 ;
  assign mem[919 ] = 5'h10 ;
  assign mem[920 ] = 5'h00 ;
  assign mem[921 ] = 5'h02 ;
  assign mem[922 ] = 5'h11 ;
  assign mem[923 ] = 5'h10 ;
  assign mem[924 ] = 5'h00 ;
  assign mem[925 ] = 5'h01 ;
  assign mem[926 ] = 5'h10 ;
  assign mem[927 ] = 5'h00 ;
  assign mem[928 ] = 5'h04 ;
  assign mem[929 ] = 5'h13 ;
  assign mem[930 ] = 5'h12 ;
  assign mem[931 ] = 5'h11 ;
  assign mem[932 ] = 5'h10 ;
  assign mem[933 ] = 5'h00 ;
  assign mem[934 ] = 5'h01 ;
  assign mem[935 ] = 5'h10 ;
  assign mem[936 ] = 5'h00 ;
  assign mem[937 ] = 5'h02 ;
  assign mem[938 ] = 5'h11 ;
  assign mem[939 ] = 5'h10 ;
  assign mem[940 ] = 5'h00 ;
  assign mem[941 ] = 5'h01 ;
  assign mem[942 ] = 5'h10 ;
  assign mem[943 ] = 5'h00 ;
  assign mem[944 ] = 5'h03 ;
  assign mem[945 ] = 5'h12 ;
  assign mem[946 ] = 5'h11 ;
  assign mem[947 ] = 5'h10 ;
  assign mem[948 ] = 5'h00 ;
  assign mem[949 ] = 5'h01 ;
  assign mem[950 ] = 5'h10 ;
  assign mem[951 ] = 5'h00 ;
  assign mem[952 ] = 5'h02 ;
  assign mem[953 ] = 5'h11 ;
  assign mem[954 ] = 5'h10 ;
  assign mem[955 ] = 5'h00 ;
  assign mem[956 ] = 5'h01 ;
  assign mem[957 ] = 5'h10 ;
  assign mem[958 ] = 5'h00 ;
  assign mem[959 ] = 5'h05 ;
  assign mem[960 ] = 5'h14 ;
  assign mem[961 ] = 5'h13 ;
  assign mem[962 ] = 5'h12 ;
  assign mem[963 ] = 5'h11 ;
  assign mem[964 ] = 5'h10 ;
  assign mem[965 ] = 5'h00 ;
  assign mem[966 ] = 5'h01 ;
  assign mem[967 ] = 5'h10 ;
  assign mem[968 ] = 5'h00 ;
  assign mem[969 ] = 5'h02 ;
  assign mem[970 ] = 5'h11 ;
  assign mem[971 ] = 5'h10 ;
  assign mem[972 ] = 5'h00 ;
  assign mem[973 ] = 5'h01 ;
  assign mem[974 ] = 5'h10 ;
  assign mem[975 ] = 5'h00 ;
  assign mem[976 ] = 5'h03 ;
  assign mem[977 ] = 5'h12 ;
  assign mem[978 ] = 5'h11 ;
  assign mem[979 ] = 5'h10 ;
  assign mem[980 ] = 5'h00 ;
  assign mem[981 ] = 5'h01 ;
  assign mem[982 ] = 5'h10 ;
  assign mem[983 ] = 5'h00 ;
  assign mem[984 ] = 5'h02 ;
  assign mem[985 ] = 5'h11 ;
  assign mem[986 ] = 5'h10 ;
  assign mem[987 ] = 5'h00 ;
  assign mem[988 ] = 5'h01 ;
  assign mem[989 ] = 5'h10 ;
  assign mem[990 ] = 5'h00 ;
  assign mem[991 ] = 5'h04 ;
  assign mem[992 ] = 5'h13 ;
  assign mem[993 ] = 5'h12 ;
  assign mem[994 ] = 5'h11 ;
  assign mem[995 ] = 5'h10 ;
  assign mem[996 ] = 5'h00 ;
  assign mem[997 ] = 5'h01 ;
  assign mem[998 ] = 5'h10 ;
  assign mem[999 ] = 5'h00 ;
  assign mem[1000] = 5'h02 ;
  assign mem[1001] = 5'h11 ;
  assign mem[1002] = 5'h10 ;
  assign mem[1003] = 5'h00 ;
  assign mem[1004] = 5'h01 ;
  assign mem[1005] = 5'h10 ;
  assign mem[1006] = 5'h00 ;
  assign mem[1007] = 5'h03 ;
  assign mem[1008] = 5'h12 ;
  assign mem[1009] = 5'h11 ;
  assign mem[1010] = 5'h10 ;
  assign mem[1011] = 5'h00 ;
  assign mem[1012] = 5'h01 ;
  assign mem[1013] = 5'h10 ;
  assign mem[1014] = 5'h00 ;
  assign mem[1015] = 5'h02 ;
  assign mem[1016] = 5'h11 ;
  assign mem[1017] = 5'h10 ;
  assign mem[1018] = 5'h00 ;
  assign mem[1019] = 5'h01 ;
  assign mem[1020] = 5'h10 ;
  assign mem[1021] = 5'h00 ;
  
  //----
  generate 
  if (RD_TYPE==0)
  begin:U_type0
    reg [$clog2(D)-1:0]addr_d1;

    always @(posedge clk)
    begin
      if((!we) & ce)
        addr_d1 <= addr;
    end

    assign rdata = mem[addr_d1];
  end
  else 
  begin:U_type1

    reg [W-1:0]rdata_int;
    always @(posedge clk)
    begin
      if((!we) & ce)
        rdata_int <= mem[addr];
    end

    assign rdata = rdata_int;
  end
  endgenerate
endmodule
